�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Pclassq0X   Sexq1X   Ageq2X   SibSpq3X   Parchq4X   Fareq5X   Embarkedq6etq7bX   n_features_in_q8KX
   n_outputs_q9KX   classes_q:h"h#K �q;h%�q<Rq=(KK�q>h)X   i8q?���q@RqA(KX   <qBNNNJ����J����K tqCb�C               qDtqEbX
   n_classes_qFKX   base_estimator_qGhX   estimators_qH]qI(h)�qJ}qK(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h8Kh9Kh:h"h#K �qLh%�qMRqN(KK�qOh)X   f8qP���qQRqR(KhBNNNJ����J����K tqSb�C              �?qTtqUbhFcnumpy.core.multiarray
scalar
qVhAC       qW�qXRqYX   max_features_qZKX   tree_q[csklearn.tree._tree
Tree
q\Kh"h#K �q]h%�q^Rq_(KK�q`hA�C       qatqbbK�qcRqd}qe(hKX
   node_countqfK�X   nodesqgh"h#K �qhh%�qiRqj(KK��qkh)X   V56ql���qmRqn(Kh-N(X
   left_childqoX   right_childqpX   featureqqX	   thresholdqrX   impurityqsX   n_node_samplesqtX   weighted_n_node_samplesqutqv}qw(hoh)X   i8qx���qyRqz(KhBNNNJ����J����K tq{bK �q|hphzK�q}hqhzK�q~hrhRK�qhshRK �q�hthzK(�q�huhRK0�q�uK8KKtq�b�B8#         @                     @zV�O6��?           �{@       +                    �?      �?t            �f@                           �?d}h��?H             \@                           �?�\��N��?             3@       
                 �|�=@��S���?             .@       	                     �?؇���X�?             @                        ȈP@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �?      �?              @                           �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                          �8@      �?             @������������������������       �                     @������������������������       �                     �?                           �?<)�%�w�?:            @W@                          �'@�LQ�1	�?             7@                          �F@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     2@       $                     �?������?+            �Q@       #                   �F@؇���X�?            �A@                            A@�E��ӭ�?             2@                           <@�8��8��?             (@������������������������       �                     @                          �>@z�G�z�?             @������������������������       �                     �?������������������������       �                     @!       "                 ��I*@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             1@%       &                 �|Y=@(N:!���?            �A@������������������������       �                     1@'       *                   @A@�<ݚ�?             2@(       )                 `fF)@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@,       ?                    �?      �?,             Q@-       .                    �?�2�o�U�?$            �K@������������������������       �                     8@/       0                    %@`՟�G��?             ?@������������������������       �                     @1       8                   �G@��}*_��?             ;@2       3                 0�"K@�<ݚ�?             2@������������������������       �                     "@4       7                     �?X�<ݚ�?             "@5       6                 03�M@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @9       :                    �?�q�q�?             "@������������������������       �                     @;       >                    �?      �?             @<       =                   @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@A       Z                   �0@�x��6�?�            �p@B       G                    �?�û��|�?             G@C       F                    '@ףp=
�?             $@D       E                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @H       M                    �?      �?             B@I       L                 P��@؇���X�?             @J       K                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @N       Q                     @ܷ��?��?             =@O       P                    #@�q�q�?             @������������������������       �                      @������������������������       �                     @R       S                    �?�nkK�?             7@������������������������       �                     @T       Y                    �?�IєX�?	             1@U       V                    @z�G�z�?             @������������������������       �                      @W       X                 ��T?@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@[       v                    �?�	{���?�            @k@\       o                    �?�ݜ����?$            �M@]       `                 �Y5@�99lMt�?            �C@^       _                 03�@�IєX�?
             1@������������������������       �                     �?������������������������       �        	             0@a       n                 �|Y>@8�A�0��?             6@b       m                    �?      �?             2@c       h                    �?     ��?             0@d       e                    �?      �?              @������������������������       �                     @f       g                    �?���Q��?             @������������������������       �                      @������������������������       �                     @i       j                   �3@      �?              @������������������������       �                      @k       l                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @p       u                    @R���Q�?             4@q       t                 0C�3@      �?             (@r       s                 ��"@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @w       �                 �?�@,_ʯ08�?a            �c@x       �                    �?��+��<�?4            �U@y       �                    �?Ћ����?1            �T@z       {                   �5@�LQ�1	�?             7@������������������������       �                     �?|       �                   @@�C��2(�?             6@}       ~                 ���@���N8�?
             5@������������������������       �                      @       �                 �|�=@$�q-�?             *@�       �                 �|=@�����H�?             "@������������������������       �                     @������������������������       �r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        %            �M@������������������������       �                     @�       �                   @E@d1<+�C�?-            @R@�       �                 �|Y=@�U�=���?)            �P@�       �                    �?r�q��?             8@�       �                 ���@@      �?             0@�       �                 ���"@��S�ۿ?             .@������������������������       �        	             (@�       �                    8@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                 @a&@      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?�Ń��̧?             E@�       �                    �? ��WV�?             :@�       �                 @3�@ �q�q�?             8@������������������������       �                     �?������������������������       �                     7@������������������������       �                      @������������������������       �                     0@�       �                 ��!@����X�?             @�       �                 @3�@r�q��?             @������������������������       �                     @�       �                   @F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KK�KK�q�hR�B
       pr@     �b@     �V@     �V@     @R@     �C@      "@      $@       @      @      @      �?      @      �?              �?      @               @               @      @      �?      @              @      �?              �?              �?      @              @      �?              P@      =@      @      4@      @       @               @      @                      2@     �N@      "@      >@      @      *@      @      &@      �?      @              @      �?              �?      @               @      @       @                      @      1@              ?@      @      1@              ,@      @       @      @       @                      @      (@              1@     �I@      1@      C@              8@      1@      ,@              @      1@      $@      ,@      @      "@              @      @      @      @              @      @               @              @      @              @      @      �?       @      �?       @                      �?      �?                      *@     �i@     �M@      <@      2@      �?      "@      �?      @              @      �?                      @      ;@      "@      �?      @      �?      �?              �?      �?                      @      :@      @      @       @               @      @              6@      �?      @              0@      �?      @      �?       @               @      �?       @                      �?      (@              f@     �D@      ?@      <@      ,@      9@      �?      0@      �?                      0@      *@      "@      "@      "@      @      "@       @      @              @       @      @       @                      @      @      @               @      @      �?      @                      �?       @              @              1@      @      "@      @       @      @       @                      @      @               @             @b@      *@     �T@      @     �S@      @      4@      @              �?      4@       @      4@      �?       @              (@      �?       @      �?      @              @      �?      @                      �?     �M@              @             �O@      $@     �N@      @      4@      @      ,@       @      ,@      �?      (@               @      �?       @                      �?              �?      @       @               @      @             �D@      �?      9@      �?      7@      �?              �?      7@               @              0@               @      @      �?      @              @      �?       @      �?                       @      �?        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfK�hgh"h#K �q�h%�q�Rq�(KK��q�hn�B�%                             #@^H���+�?           �{@                           �?R�}e�.�?             :@������������������������       �        
             3@������������������������       �                     @       N                     @Ƈ���3�?            z@                           �?X�����?o             f@       
                   �'@ �.�?Ƞ?#             N@       	                   �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        !            �L@                           -@&d���?L             ]@������������������������       �                      @       +                 ��D:@L�}�:G�?K            �\@                           �?�:pΈ��?#             I@                           �?      �?             @                        �|Y:@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?       *                    �?�q��/��?              G@       )                    �?,���i�?            �D@       &                   �D@      �?             D@                           @�KM�]�?             C@������������������������       �                     @                            �?��� ��?             ?@������������������������       �                      @                           &@\-��p�?             =@                          �5@�q�q�?             @������������������������       �                      @������������������������       �                     @        !                   �(@���}<S�?             7@������������������������       �                     @"       #                 �|�<@�KM�]�?             3@������������������������       �                     $@$       %                   �@@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @'       (                 `f�)@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @,       I                   �I@     ��?(             P@-       <                   �@@(옄��?             G@.       5                 �|�<@z�G�z�?             9@/       0                   �8@@4և���?             ,@������������������������       �                      @1       4                    �?r�q��?             @2       3                 ��3Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @6       ;                 �|Y>@���|���?             &@7       8                    �?X�<ݚ�?             "@������������������������       �                     @9       :                   �D@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @=       H                   �G@���N8�?             5@>       ?                    �?X�Cc�?             ,@������������������������       �                     @@       G                    �?X�<ݚ�?             "@A       F                     �?����X�?             @B       E                    F@�q�q�?             @C       D                  x#J@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @J       K                 ȈP@�X�<ݺ?             2@������������������������       �                     *@L       M                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @O       �                    �?����?�            @n@P       �                   @@@�>:���?�            `l@Q       �                 0��F@���]�3�?t             g@R       �                    �?ƆQ����?r            �f@S       X                   �0@�0���?f            �d@T       U                    '@��
ц��?             *@������������������������       �                     �?V       W                    �?      �?             (@������������������������       �                     @������������������������       �                     @Y       �                   �>@>A�F<�?_             c@Z       i                    �?��H�&p�?]            �b@[       `                    �?�lg����?            �E@\       _                 `fV&@z�G�z�?
             .@]       ^                 �|�7@$�q-�?	             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                      @a       h                 �|Y=@؇���X�?             <@b       g                 �Y�@���Q��?             $@c       f                    �?؇���X�?             @d       e                   @8@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     2@j       �                    �?0��_��?A            �Z@k       l                   �5@ 	��p�?6            �U@������������������������       �                     7@m       �                 ���"@     ��?'             P@n       s                    �? 	��p�?"             M@o       r                  sW@      �?             @p       q                   �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?t       u                   �7@�X�<ݺ?             K@������������������������       �                     .@v       y                 ���@$�q-�?            �C@w       x                 �|�:@      �?             @������������������������       �                      @������������������������       �                      @z                        �?$@��?^�k�?            �A@{       |                 pf�@�C��2(�?             &@������������������������       �                      @}       ~                 �|Y=@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    (@���Q��?             @�       �                   �:@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �!@���y4F�?             3@�       �                    �?���Q��?             $@������������������������       �                     �?�       �                    5@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                 ��� @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 ��*@X�<ݚ�?             2@�       �                 �|Y<@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                 `v�6@"pc�
�?	             &@�       �                    5@����X�?             @������������������������       �                     @�       �                    @      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?@4և���?             E@�       �                   �E@ >�֕�?            �A@������������������������       �                     9@�       �                   @F@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                      @�       �                   @A@z�G�z�?             @������������������������       �                      @�       �                 0336@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             .@q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hR�B�
        r@     �c@      @      3@              3@      @             �q@      a@     �U@     �V@      �?     �M@      �?       @               @      �?                     �L@     @U@      ?@               @     @U@      =@     �E@      @       @       @      �?       @      �?                       @      �?             �D@      @      B@      @     �A@      @      A@      @      @              ;@      @       @              9@      @      @       @               @      @              5@       @      @              1@       @      $@              @       @               @      @              �?      �?      �?                      �?      �?              @              E@      6@      9@      5@      4@      @      *@      �?       @              @      �?      �?      �?              �?      �?              @              @      @      @      @      @              �?      @              @      �?               @              @      0@      @      "@              @      @      @      @       @      @       @      @       @      @                       @      �?              �?                       @              @      1@      �?      *@              @      �?              �?      @             `h@     �G@     �f@     �G@     �a@      F@     �a@      E@     ``@      A@      @      @      �?              @      @              @      @              _@      <@     �^@      :@      ;@      0@      @      (@      �?      (@      �?                      (@       @              8@      @      @      @      @      �?      @      �?              �?      @              @                      @      2@              X@      $@     @T@      @      7@              M@      @      K@      @      @      �?       @      �?              �?       @              �?             �I@      @      .@              B@      @       @       @               @       @              A@      �?      $@      �?       @               @      �?       @                      �?      8@              @       @      �?              @       @      �?       @      �?                       @       @              .@      @      @      @              �?      @      @              @      @              "@              �?       @      �?                       @      $@       @      �?      @              @      �?              "@       @      @       @      @               @       @      �?       @               @      �?              �?              @                       @     �C@      @     �@@       @      9@               @       @               @       @              @      �?       @              @      �?       @               @      �?              �?       @              .@        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfK�hgh"h#K �q�h%�q�Rq�(KK��q�hn�B�%         *                    �?�Gi����?           �{@       )                    �?��9܂�?7            @V@       
                    �?j���� �?6            @U@                            @�C��2(�?            �@@������������������������       �                     :@                          �+@և���X�?             @������������������������       �                      @       	                    �?���Q��?             @������������������������       �                     @������������������������       �                      @                            �?�n_Y�K�?              J@                          �8@և���X�?             5@������������������������       �                      @                           �?�	j*D�?
             *@                        �D@E@�q�q�?             @������������������������       �                      @                           �?      �?             @������������������������       �                      @������������������������       �                      @                        ���X@����X�?             @������������������������       �                     @������������������������       �                      @                          �5@f���M�?             ?@������������������������       �                     @                            @z�G�z�?             9@                        hf�2@�q�q�?             @������������������������       �                     �?������������������������       �                      @       $                   @@"pc�
�?             6@                        ���@�X�<ݺ?
             2@������������������������       �                      @        !                 �|=@ףp=
�?             $@������������������������       �                     @"       #                 �|�=@r�q��?             @������������������������       �z�G�z�?             @������������������������       �                     �?%       (                 ��*@      �?             @&       '                 �|Y=@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       X                     @"` Y��?�            0v@,       /                    �?�C�gOS�?[             c@-       .                   �'@0�)AU��?%            �L@������������������������       �                     �?������������������������       �        $             L@0       G                     �?�q�q��?6             X@1       F                    @v ��?            �E@2       E                   @J@��6���?             E@3       4                   �9@�!���?             A@������������������������       �                     @5       D                    �?�>4և��?             <@6       =                   �@@�q�q�?             8@7       8                 0�D@X�<ݚ�?             "@������������������������       �                     @9       :                    �?z�G�z�?             @������������������������       �                     @;       <                    9@      �?              @������������������������       �                     �?������������������������       �                     �?>       ?                    �?��S�ۿ?             .@������������������������       �                     (@@       A                 0�nL@�q�q�?             @������������������������       �                     �?B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?H       U                    �?�#ʆA��?            �J@I       T                    �?R���Q�?             D@J       K                 `f�)@���!pc�?            �@@������������������������       �                     &@L       M                 �|Y<@8�A�0��?	             6@������������������������       �                     $@N       S                   @D@      �?             (@O       R                   �3@      �?             @P       Q                   �A@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @V       W                    &@��
ц��?             *@������������������������       �                     @������������������������       �                     @Y       �                    �?.p����?�            @i@Z       q                   �;@�G��l��?#             E@[       h                    �?���|���?             6@\       g                   �6@؇���X�?             ,@]       f                    �?�<ݚ�?	             "@^       _                    1@����X�?             @������������������������       �                      @`       a                 ���@���Q��?             @������������������������       �                     �?b       c                   �5@      �?             @������������������������       �                      @d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @i       n                    @      �?              @j       m                    �?r�q��?             @k       l                 �!@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @o       p                 ��T?@      �?              @������������������������       �                     �?������������������������       �                     �?r                           B@�z�G��?             4@s       ~                   �@@      �?             0@t       }                    �?����X�?             ,@u       v                 �|�<@      �?              @������������������������       �                     �?w       |                 �|Y>@և���X�?             @x       y                 ���@      �?             @������������������������       �                     �?z       {                 `f�@���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?ףp=
�?_             d@������������������������       �                     =@�       �                    @��ϻ�r�?Q            ``@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 @3�@     ��?O             `@������������������������       �                     @�       �                    �?h�N?���?N            @_@�       �                 �T)D@@��xQ�?F            �\@�       �                    �?��X��?E             \@�       �                    �?��-#���?A            �Z@�       �                 pF� @�c:��?9             W@�       �                   �E@��IF�E�?-            �P@�       �                 �?�@ 	��p�?(             M@�       �                    9@��?^�k�?            �A@�       �                   �7@      �?             0@������������������������       �        	             ,@�       �                   �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@�       �                 @3�@�LQ�1	�?             7@������������������������       �                     �?�       �                   �4@�C��2(�?             6@�       �                   �1@�q�q�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     0@�       �                 pff@      �?              @������������������������       �                     @�       �                 @3�@      �?             @������������������������       �                      @�       �                   @F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     :@�       �                 P�@؇���X�?             ,@������������������������       �                     @�       �                 ��y'@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     &@q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hR�B�
       �p@     �f@     �C@      I@     �A@      I@      @      >@              :@      @      @               @      @       @      @                       @      @@      4@      (@      "@       @              @      "@       @      @               @       @       @       @                       @       @      @              @       @              4@      &@              @      4@      @       @      �?              �?       @              2@      @      1@      �?       @              "@      �?      @              @      �?      @      �?      �?              �?      @      �?       @               @      �?                      �?      @              l@     @`@     �M@     �W@      �?      L@      �?                      L@      M@      C@      4@      7@      3@      7@      &@      7@      @              @      7@      @      3@      @      @              @      @      �?      @              �?      �?      �?                      �?      �?      ,@              (@      �?       @              �?      �?      �?      �?                      �?              @       @              �?              C@      .@      ?@      "@      8@      "@      &@              *@      "@      $@              @      "@      @      @       @      @              @       @              �?                      @      @              @      @              @      @             �d@      B@      6@      4@       @      ,@       @      (@       @      @       @      @               @       @      @      �?              �?      @               @      �?      �?              �?      �?                       @              @      @       @      @      �?       @      �?              �?       @              @              �?      �?      �?                      �?      ,@      @      $@      @      $@      @      @      @      �?              @      @      @      @              �?      @       @       @       @      �?                      �?      @                       @      @              b@      0@      =@             �\@      0@      �?       @               @      �?             �\@      ,@              @     �\@      &@     �Y@      &@     �Y@      "@     @X@      "@     @U@      @     �M@      @      K@      @      A@      �?      .@      �?      ,@              �?      �?              �?      �?              3@              4@      @              �?      4@       @      @       @      @              �?       @      0@              @      @      @              �?      @               @      �?      �?      �?                      �?      :@              (@       @      @              @       @               @      @              @                       @      &@        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       qՆq�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfK�hgh"h#K �q�h%�q�Rq�(KK��q�hn�B�)         t                 Ь�9@Z�.!c��?           �{@                          �0@����;�?�             q@       
                 ��*4@�+e�X�?             9@       	                 ��.#@؇���X�?             5@                        ��@���!pc�?             &@������������������������       �                     @                        pf�@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �        	             $@                            @      �?             @������������������������       �                     �?������������������������       �                     @       a                   �?@*��r��?�            �n@       J                 `f�%@���N8�?}            �g@       '                    �?z�G�z�?Z            �`@                          �6@j���� �?             A@������������������������       �                     @                          �<@f���M�?             ?@������������������������       �                     @                           �?
j*D>�?             :@                        pF @�	j*D�?	             *@                           �?ףp=
�?             $@������������������������       �                     �?                        ���@�����H�?             "@������������������������       �                     �?                        �&B@      �?              @������������������������       �؇���X�?             @������������������������       �                     �?������������������������       �                     @       $                 03s@8�Z$���?             *@        #                    �?�C��2(�?
             &@!       "                 ���@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@%       &                 �|Y=@      �?              @������������������������       �                     �?������������������������       �                     �?(       5                 �Yu@�_�s���?A            @Y@)       *                     @��s����?             E@������������������������       �                     @+       4                   �8@x�����?            �C@,       -                    �?���|���?             6@������������������������       �                     @.       3                    �?      �?	             0@/       2                 ���@8�Z$���?             *@0       1                   �5@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @������������������������       �        
             1@6       G                   �>@�U�:��?'            �M@7       8                     @�h����?%             L@������������������������       �                     @9       @                   �<@ �h�7W�?#            �J@:       ;                    �?��?^�k�?            �A@������������������������       �                     "@<       =                    �? ��WV�?             :@������������������������       �                     6@>       ?                    8@      �?             @������������������������       �                     �?������������������������       �                     @A       B                 ��) @�����H�?             2@������������������������       �        	             .@C       D                 pf� @�q�q�?             @������������������������       �                     �?E       F                 ��)"@      �?              @������������������������       �                     �?������������������������       �                     �?H       I                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @K       V                     @�q�q�?#             K@L       M                    �?և���X�?             <@������������������������       �                      @N       O                   �(@z�G�z�?             4@������������������������       �                     @P       S                    �?      �?             0@Q       R                 `��,@z�G�z�?             @������������������������       �                     �?������������������������       �                     @T       U                 �|�<@���!pc�?             &@������������������������       �                      @������������������������       �                     @W       X                 ��*@�θ�?             :@������������������������       �                     @Y       Z                 �=/@�C��2(�?             6@������������������������       �                     @[       `                    �?�r����?
             .@\       ]                 �2@�q�q�?             @������������������������       �                     �?^       _                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@b       s                    �?��ϭ�*�?$             M@c       d                    �?�Ra����?             F@������������������������       �                     "@e       l                    �?؇���X�?            �A@f       k                    �?�q�q�?             "@g       j                     @և���X�?             @h       i                   @H@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @m       n                 �?�@$�q-�?             :@������������������������       �                     (@o       p                   @F@؇���X�?	             ,@������������������������       �                     &@q       r                 ��!@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             ,@u       �                 �U�R@�����?l            �e@v       �                    �?��S���?M             ^@w       �                     @�q�����?>             Y@x       �                   �J@`՟�G��?9            @W@y       �                    �?$��m��?0            �S@z       {                 ���=@      �?             $@������������������������       �                     �?|       �                   �H@X�<ݚ�?             "@}       ~                     �?և���X�?             @������������������������       �                     @       �                   �7@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�!���?(             Q@�       �                     �?��?^�k�?            �A@������������������������       �                     *@�       �                    �?���7�?
             6@�       �                   @B@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�       �                   �>@���|���?            �@@�       �                    �?���Q��?             .@�       �                     �?"pc�
�?	             &@�       �                 ��$:@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?������������������������       �                     @�       �                    �?r�q��?             2@������������������������       �                      @�       �                   @B@�z�G��?             $@������������������������       �                     @�       �                 0�nL@և���X�?             @�       �                  x#J@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             .@�       �                 0�H@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                 ��p@@z�G�z�?             4@�       �                    �?���|���?             &@������������������������       �                      @�       �                    @X�<ݚ�?             "@������������������������       �                     @�       �                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                 `fmj@R�}e�.�?             J@�       �                    �?&^�)b�?            �E@������������������������       �                     <@�       �                    �?��S���?	             .@�       �                   @B@���!pc�?             &@������������������������       �                     @�       �                    L@      �?             @�       �                   �I@���Q��?             @�       �                 ���X@�q�q�?             @������������������������       �                     �?�       �                   �H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             "@������������������������       �                      @�       �                    �?؇���X�?             @�       �                 X�l@@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hR�B�       �q@     `d@     `i@     @Q@      @      3@      @      2@      @       @              @      @       @       @              �?       @              $@      @      �?              �?      @             �h@      I@      b@     �F@      [@      ;@      4@      ,@              @      4@      &@      @              .@      &@      @      "@      �?      "@              �?      �?       @              �?      �?      @      �?      @              �?      @              &@       @      $@      �?      �?      �?      �?                      �?      "@              �?      �?              �?      �?              V@      *@      A@       @      @              ?@       @      ,@       @              @      ,@       @      &@       @      �?       @      �?                       @      $@              @              1@              K@      @     �J@      @      @              I@      @      A@      �?      "@              9@      �?      6@              @      �?              �?      @              0@       @      .@              �?       @              �?      �?      �?      �?                      �?      �?       @      �?                       @      B@      2@      0@      (@               @      0@      @      @              (@      @      @      �?              �?      @               @      @       @                      @      4@      @              @      4@       @      @              *@       @      �?       @              �?      �?      �?              �?      �?              (@             �J@      @     �C@      @      "@              >@      @      @      @      @      @      @      @              @      @              �?               @              8@       @      (@              (@       @      &@              �?       @               @      �?              ,@             �S@     �W@      P@      L@      H@      J@      E@     �I@      ;@     �I@      @      @              �?      @      @      @      @              @      @      �?              �?      @               @              6@      G@      �?      A@              *@      �?      5@      �?      @              @      �?                      .@      5@      (@      @      "@       @      "@      �?      "@      �?                      "@      �?              @              .@      @       @              @      @      @              @      @      �?      @      �?                      @      @              .@              @      �?      @                      �?      0@      @      @      @       @              @      @      @              �?      @      �?                      @      "@              ,@      C@       @     �A@              <@       @      @       @      @      @              @      @      @       @      �?       @              �?      �?      �?      �?                      �?       @                      �?              @      @      @               @      @      �?      @      �?      @                      �?       @        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}r   (hKhfK�hgh"h#K �r  h%�r  Rr  (KK��r  hn�B$         >                     @^H���+�?           �{@                          �1@��hX���?r            �f@������������������������       �                     1@                           �?�W1���?g            �d@                          �'@     p�?,             P@                          �F@      �?             @������������������������       �                     �?������������������������       �                     @	       
                   �E@(;L]n�?*             N@������������������������       �        "            �G@                         x�C@8�Z$���?             *@                           �?���Q��?             @                            �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @       '                    A@z�G�z�?;             Y@       &                 ���=@l�b�G��?#            �L@                           4@��� ��?             ?@                           &@      �?              @������������������������       �                     �?������������������������       �                     �?                            �?ܷ��?��?             =@                        ���;@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        `fF)@$�q-�?             :@������������������������       �                     *@       %                    �?8�Z$���?             *@       "                    �?�<ݚ�?             "@        !                 ���,@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                   �=@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     :@(       )                    B@�lg����?            �E@������������������������       �                     @*       =                    �?����>�?            �B@+       <                 ���S@�E��ӭ�?             B@,       ;                   @M@�'�`d�?            �@@-       :                    �?�q�q�?             5@.       /                 ��:@j���� �?
             1@������������������������       �                     @0       9                   �K@��
ц��?             *@1       8                     �?�eP*L��?             &@2       7                   �J@      �?             $@3       4                 03�C@����X�?             @������������������������       �                     @5       6                  x#J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     (@������������������������       �                     @������������������������       �                     �??       @                    �?ҹ��!��?�            pp@������������������������       �                     @A       �                    �?��j����?�            @p@B       C                     @� ��Z�?�            �k@������������������������       �                     @D       �                 �T�I@Ƶ�pD�?�             k@E       �                    �?H芦��?�            �j@F       U                    �?^$T�|��?y             h@G       P                 �|Y=@�q����?            �J@H       O                 �&�)@�G��l��?
             5@I       N                 �Y�@������?             .@J       M                   �5@�q�q�?             @K       L                 �Y�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     @Q       T                    �?     ��?             @@R       S                 ���@����X�?             @������������������������       �                      @������������������������       ����Q��?             @������������������������       �                     9@V       c                    �?������?[            �a@W       ^                    8@�q�q�?             8@X       ]                   �4@�	j*D�?             *@Y       \                   �3@և���X�?             @Z       [                    0@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @_       b                    �?�C��2(�?             &@`       a                 ��� @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @d       �                    �?��Õty�?M             ]@e       �                   @C@\�t��Y�?D            �Y@f       i                   �0@|)����?:            �V@g       h                 pf�@      �?             @������������������������       �                      @������������������������       �      �?              @j       s                   �7@����?7            �U@k       r                   �3@г�wY;�?             A@l       m                   �2@�C��2(�?
             &@������������������������       �                     @n       o                 �?�@      �?              @������������������������       �                     @p       q                 `�8"@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     7@t       u                  ��	@���C��?             �J@������������������������       �                     �?v       �                 �|�=@4��?�?             J@w       ~                 �?$@,���i�?            �D@x       y                   �8@�θ�?             *@������������������������       �                     �?z       {                 �|Y=@r�q��?             (@������������������������       �                     @|       }                 ��@      �?              @������������������������       �                     @������������������������       �                      @       �                 ��)"@@4և���?             <@������������������������       �                     3@�       �                   �<@�<ݚ�?             "@������������������������       �                     @�       �                 �|Y=@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     &@�       �                 pff@�q�q�?
             (@������������������������       �                     @�       �                    G@և���X�?             @�       �                 pf� @�q�q�?             @�       �                   @F@z�G�z�?             @�       �                 @3�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    5@$�q-�?	             *@������������������������       �                     �?������������������������       �                     (@�       �                    @�eP*L��?             6@�       �                    �?      �?             0@�       �                 �|Y<@X�<ݚ�?             "@�       �                    @����X�?             @�       �                 ��*@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?����X�?             @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                    �B@r  tr  bh�h"h#K �r  h%�r  Rr	  (KK�KK�r
  hR�BP
        r@     �c@     @U@      X@              1@     @U@     �S@      @     �M@      @      �?              �?      @               @      M@             �G@       @      &@       @      @       @       @               @       @                      �?               @      T@      4@     �J@      @      ;@      @      �?      �?              �?      �?              :@      @       @      �?       @                      �?      8@       @      *@              &@       @      @       @       @      �?              �?       @              @      �?      @                      �?      @              :@              ;@      0@              @      ;@      $@      :@      $@      :@      @      ,@      @      $@      @      @              @      @      @      @      @      @       @      @              @       @      �?       @                      �?      @              �?                       @      @              (@                      @      �?             `i@      N@              @     `i@     �L@     �d@     �L@              @     �d@     �I@     �d@     �H@     @c@     �C@     �B@      0@      $@      &@      @      &@      @       @      �?       @      �?                       @      @                      "@      @              ;@      @       @      @               @       @      @      9@             @]@      7@      ,@      $@      @      "@      @      @      �?      @      �?                      @      @                      @      $@      �?      @      �?      @                      �?      @             �Y@      *@     �V@      (@     �T@       @      @      �?       @              �?      �?      T@      @     �@@      �?      $@      �?      @              @      �?      @               @      �?              �?       @              7@             �G@      @              �?     �G@      @      B@      @      $@      @              �?      $@       @      @              @       @      @                       @      :@       @      3@              @       @      @              @       @               @      @              &@               @      @      @              @      @       @      @      �?      @      �?       @               @      �?                       @      �?              �?              (@      �?              �?      (@              (@      $@      @      $@      @      @       @      @       @      @              @       @                      �?       @               @      @              @       @       @               @       @              @                       @     �B@        r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfK�hgh"h#K �r!  h%�r"  Rr#  (KK��r$  hn�BX)         6                    �?b��H���?           �{@       1                 ��H@节>t�?Y            �b@       "                    �?�2�o�U�?B            �[@                          �;@@�0�!��?'             Q@                           �?�IєX�?             A@                           8@HP�s��?             9@                        P�>,@���N8�?             5@������������������������       �        	             1@	       
                     @      �?             @������������������������       �                     @������������������������       �                     �?                         @$@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@       !                   �'@�t����?             A@                           �?      �?             4@                           �?"pc�
�?             &@������������������������       �                     �?                        pF @z�G�z�?             $@                        ���@�����H�?             "@������������������������       �                     �?                        �&B@      �?              @������������������������       �؇���X�?             @������������������������       �                     �?������������������������       �                     �?                        �|�?@�����H�?             "@������������������������       �                     @                        `f$@z�G�z�?             @������������������������       �                     @                           �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@#       $                     @�G��l��?             E@������������������������       �                     0@%       0                    @8�Z$���?             :@&       /                    �?"pc�
�?             6@'       (                   �$@���Q��?             $@������������������������       �                      @)       *                 �|Y9@      �?              @������������������������       �                     @+       ,                  S�-@���Q��?             @������������������������       �                     �?-       .                 �|�>@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     (@������������������������       �                     @2       5                 �|�=@�7��?            �C@3       4                     @�t����?	             1@������������������������       �                     .@������������������������       �                      @������������������������       �                     6@7       b                     �?�d���?�            pr@8       I                    �? 1_#�?%            �M@9       :                   �8@�\��N��?             3@������������������������       �                     @;       B                    �?     ��?	             0@<       A                    �?      �?              @=       @                   �O@և���X�?             @>       ?                 `fp`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?C       H                 ���X@      �?              @D       E                 ���S@r�q��?             @������������������������       �                     @F       G                 ��hU@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @J       _                    �?R���Q�?             D@K       ^                    �?b�h�d.�?            �A@L       M                   @A@��hJ,�?             A@������������������������       �                     $@N       ]                    �?�q�q�?             8@O       V                 `f�;@�GN�z�?             6@P       U                    J@X�<ݚ�?             "@Q       T                   @E@�q�q�?             @R       S                 ��I*@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @W       X                    �?$�q-�?             *@������������������������       �                     $@Y       Z                  x#J@�q�q�?             @������������������������       �                     �?[       \                    F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?`       a                    @���Q��?             @������������������������       �                     @������������������������       �                      @c       f                    @p/3�d��?�            �m@d       e                   �;@      �?             0@������������������������       �                     (@������������������������       �                     @g       ~                 �?�@ףp=
�?�            �k@h       q                    �? �#�Ѵ�?7            �U@i       j                   �5@�θ�?	             *@������������������������       �                     �?k       p                 �|�=@r�q��?             (@l       m                 ���@�<ݚ�?             "@������������������������       �                     @n       o                 �|�:@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     @r       s                 �|Y=@ �й���?.            @R@������������������������       �                     ;@t       u                     @��<b�ƥ?             G@������������������������       �                      @v       w                    �?`���i��?             F@������������������������       �                     3@x       }                  sW@`2U0*��?             9@y       |                 �|�?@�����H�?             "@z       {                 pf�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@       �                 @3�@��v����?]            �`@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �4@     ��?Y             `@�       �                     @d}h���?             <@�       �                    �?�����?             3@�       �                     @      �?             0@�       �                   �2@r�q��?             @������������������������       �                     @�       �                   �'@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 pf� @�z�G��?             $@�       �                   �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    )@�q�q�?             @������������������������       �                     �?�       �                 ��1@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �?HP�s��?E             Y@�       �                   �9@����X�?             @������������������������       �                      @�       �                 @Q,@���Q��?             @������������������������       �                     �?�       �                     @      �?             @������������������������       �                     �?�       �                   �:@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?`Jj��??            @W@������������������������       �                     �?�       �                 0�_F@���.�6�?>             W@�       �                 ��+@��`qM|�?7            �T@�       �                     @Hm_!'1�?"            �H@�       �                   �@@�����H�?             2@������������������������       �                     &@�       �                 `f�)@����X�?             @������������������������       �                     @�       �                   �A@      �?             @������������������������       �                     �?�       �                   @D@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �<@`Jj��?             ?@������������������������       �        	             .@�       �                 ��) @      �?             0@������������������������       �                     *@�       �                 X��@@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     A@�       �                    �?�<ݚ�?             "@�       �                   �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KK�KK�r*  hR�B�       pq@     �d@      B@     @\@      A@      S@      (@      L@       @      @@       @      7@      �?      4@              1@      �?      @              @      �?              �?      @      �?                      @              "@      $@      8@      $@      $@       @      "@              �?       @       @      �?       @              �?      �?      @      �?      @              �?      �?               @      �?      @              @      �?      @              �?      �?              �?      �?                      ,@      6@      4@              0@      6@      @      2@      @      @      @               @      @       @      @              @       @      �?               @       @               @       @              (@              @               @     �B@       @      .@              .@       @                      6@     `n@      J@     �D@      2@      $@      "@      @              @      "@      @      @      @      @      �?      @              @      �?               @              �?              @      @      �?      @              @      �?       @      �?                       @       @              ?@      "@      =@      @      =@      @      $@              3@      @      1@      @      @      @       @      @       @      �?       @                      �?              @      @              (@      �?      $@               @      �?      �?              �?      �?              �?      �?               @                      �?       @      @              @       @             @i@      A@      @      (@              (@      @             �h@      6@     �T@      @      $@      @              �?      $@       @      @       @      @              @       @       @              �?       @      @              R@      �?      ;@             �F@      �?       @             �E@      �?      3@              8@      �?       @      �?       @      �?       @                      �?      @              0@              ]@      2@       @      @              @       @             �\@      ,@      6@      @      *@      @      (@      @      @      �?      @               @      �?              �?       @              @      @      �?       @      �?                       @      @      �?      @                      �?      �?       @              �?      �?      �?              �?      �?              "@              W@       @      @       @       @              @       @              �?      @      �?      �?               @      �?              �?       @             �U@      @      �?             �U@      @     �S@      @     �F@      @      0@       @      &@              @       @      @               @       @              �?       @      �?       @                      �?      =@       @      .@              ,@       @      *@              �?       @               @      �?              A@              @       @      �?       @      �?                       @      @        r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfK�hgh"h#K �rA  h%�rB  RrC  (KKŅrD  hn�B+         F                    �?�K�n���?           �{@       A                 ��H@z�G�z�?d             d@       @                    @���?��?J            @[@       '                 `f�%@�T`�[k�?G            �Z@                           �?�q�q�?             E@                        03�@�KM�]�?             3@������������������������       �                     �?       	                 �|�9@�X�<ݺ?             2@������������������������       �                     @
                           �?@4և���?	             ,@������������������������       �                     @                        ���@�C��2(�?             &@������������������������       �                     @                        �&B@      �?              @������������������������       �r�q��?             @������������������������       �                      @                        �&B@
;&����?             7@                        ���@z�G�z�?             @������������������������       �                      @                          �7@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         Ь�#@b�2�tk�?             2@                        `�("@      �?             (@                          �9@      �?             @                        xF� @      �?             @                          �0@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @!       &                 pF%@�q�q�?             @"       #                 �yW$@z�G�z�?             @������������������������       �                     �?$       %                   �F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?(       )                    !@     ��?+             P@������������������������       �        
             ,@*       +                    -@z�G�z�?!             I@������������������������       �                      @,       =                     @r�q��?             H@-       <                    �?������?            �D@.       7                     @�J�4�?             9@/       0                    �?�C��2(�?             6@������������������������       �                     @1       2                    E@�����H�?             2@������������������������       �                     &@3       4                     �?����X�?             @������������������������       �                     @5       6                   @F@�q�q�?             @������������������������       �                      @������������������������       �                     �?8       9                 �|�;@�q�q�?             @������������������������       �                     �?:       ;                  S�-@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@>       ?                 �|�=@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @B       C                    �?���J��?            �I@������������������������       �                    �B@D       E                    @@4և���?             ,@������������������������       �                     *@������������������������       �                     �?G       j                    �?�w��.F�?�            �q@H       i                    �?      �?#             H@I       `                 ��d5@�*/�8V�?"            �G@J       M                     @��H�}�?             9@K       L                 ���,@      �?              @������������������������       �                     �?������������������������       �                     �?N       _                    �?�LQ�1	�?             7@O       T                   @;@      �?             4@P       Q                 xF*@�q�q�?             @������������������������       �                     �?R       S                   �2@      �?              @������������������������       �                     �?������������������������       �                     �?U       ^                 �|�=@@�0�!��?             1@V       W                   �<@      �?             (@������������������������       �                     @X       Y                 ���@�q�q�?             "@������������������������       �                     @Z       [                 �|Y=@���Q��?             @������������������������       �                     �?\       ]                   @@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @a       b                    A@��2(&�?             6@������������������������       �                     &@c       f                    �?���!pc�?             &@d       e                   �O@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @g       h                 ڪ�q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?k       p                    $@��lJ���?�            �m@l       m                     @��S���?	             .@������������������������       �                     @n       o                 03�6@���!pc�?             &@������������������������       �                     @������������������������       �                      @q       �                  x#J@�;��?�            �k@r       �                    �?ДX��?�            �i@s       �                 ��$:@p�/E�f�?v            �g@t       �                   �G@h7�R�
�?g            �d@u       �                    E@4��?�?a            �c@v       �                 pF� @�ma�H��?^             c@w       �                 �|�=@d۬����?:            @W@x       y                     @v���a�?0            @R@������������������������       �                     @z       �                 �?�@�� =[�?,             Q@{       �                 �?$@H�ՠ&��?#             K@|       �                    �?�'�`d�?            �@@}       �                 �|Y=@8�Z$���?	             *@~                         ��@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                 ���@      �?             4@������������������������       �                     @�       �                   @6@     ��?
             0@������������������������       �                     @�       �                    9@X�<ݚ�?             "@������������������������       �                      @�       �                 ��@և���X�?             @������������������������       �                     �?�       �                 �|Y=@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     5@�       �                    �?����X�?	             ,@�       �                    4@z�G�z�?             $@�       �                   �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        
             4@�       �                     @(;L]n�?$             N@�       �                    �?`Jj��?             ?@�       �                 �|Y=@@4և���?             <@������������������������       �        	             1@�       �                     �?"pc�
�?             &@������������������������       �                      @�       �                 �|Y?@�<ݚ�?             "@������������������������       �                     �?�       �                   @A@      �?              @�       �                   �@@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     =@�       �                 ���@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                    �?���!pc�?             6@�       �                   �J@�q�q�?             2@�       �                   �@@�eP*L��?	             &@�       �                 �|Y>@�q�q�?             @�       �                   �>@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                 03C@@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     0@�       �                    @��.k���?             1@�       �                     �?     ��?
             0@�       �                    �?      �?              @�       �                    �?����X�?             @�       �                    9@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KK�KK�rJ  hR�BP       pp@     �f@      <@     �`@      ;@     �T@      8@     �T@      ,@      <@       @      1@      �?              �?      1@              @      �?      *@              @      �?      $@              @      �?      @      �?      @               @      (@      &@      �?      @               @      �?       @               @      �?              &@      @      "@      @      @      @      @      �?      �?      �?      �?                      �?       @                       @      @               @      @      �?      @              �?      �?      @              @      �?              �?              $@      K@              ,@      $@      D@       @               @      D@      @     �B@      @      5@       @      4@              @       @      0@              &@       @      @              @       @      �?       @                      �?       @      �?      �?              �?      �?      �?                      �?              0@      @      @      @                      @      @              �?      I@             �B@      �?      *@              *@      �?             `m@     �H@      B@      (@     �A@      (@      0@      "@      �?      �?              �?      �?              .@       @      .@      @      �?       @              �?      �?      �?      �?                      �?      ,@      @      "@      @      @              @      @      @               @      @              �?       @       @      �?       @      �?              @                      @      3@      @      &@               @      @      @       @               @      @              �?      �?      �?                      �?      �?             �h@     �B@       @      @              @       @      @              @       @             �g@      >@     �f@      5@     �d@      5@     �b@      .@     �a@      .@     �a@      *@     �T@      &@      O@      &@      @             �L@      &@     �G@      @      :@      @      &@       @      @       @      @                       @       @              .@      @      @              &@      @      @              @      @               @      @      @      �?              @      @      @                      @      5@              $@      @       @       @      �?       @      �?                       @      @               @       @               @       @              4@              M@       @      =@       @      :@       @      1@              "@       @       @              @       @              �?      @      �?       @      �?       @                      �?      @              @              =@              �?       @      �?                       @      $@              0@      @      (@      @      @      @      @       @       @       @               @       @               @              �?      @              @      �?              @              @              0@               @      "@      @      "@       @      @       @      @       @      @       @                      @              �?              �?      @      @              @      @              �?        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfK�hgh"h#K �ra  h%�rb  Rrc  (KKՅrd  hn�B�.         R                     @�{S�~��?#           �{@       /                     �?���>4��?y            �h@                         x#J@Jܤm6�?A            �Y@                           �?*O���?             B@                          @M@^������?            �A@                           �?և���X�?             <@������������������������       �                     @                          �G@�q�q�?             8@	                           �?      �?             4@
                          �B@�E��ӭ�?             2@                          �>@�q�q�?             (@                           A@      �?              @                          �1@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @                           �?      �?             @������������������������       �                     �?                          �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       $                 �|Y>@:ɨ��?&            �P@                          �2@�'�=z��?            �@@������������������������       �                     @       #                 `fmj@�n_Y�K�?             :@                         ���M@X�<ݚ�?
             2@������������������������       �                      @!       "                    �?      �?	             0@������������������������       �                     $@������������������������       �                     @������������������������       �                      @%       ,                    �?<���D�?            �@@&       '                    �? �q�q�?             8@������������������������       �        
             0@(       )                    F@      �?              @������������������������       �                     @*       +                 8�<Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @-       .                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @0       1                    '@z�J��?8            �W@������������������������       �                     "@2       E                    �?,�|%�v�?3            @U@3       4                    �?��.k���?            �I@������������������������       �                     @5       6                    �?z�J��?            �G@������������������������       �        	             .@7       D                   �3@      �?             @@8       C                   @D@�LQ�1	�?             7@9       >                 `fF)@����X�?             5@:       =                    5@�C��2(�?             &@;       <                    &@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@?       @                 �|�:@      �?             $@������������������������       �                     @A       B                   �A@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     "@F       Q                    @�t����?             A@G       N                   �8@���!pc�?            �@@H       M                    �?X�<ݚ�?             "@I       J                    �?r�q��?             @������������������������       �                      @K       L                   �4@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @O       P                    �?r�q��?             8@������������������������       �                     @������������������������       �        
             4@������������������������       �                     �?S       h                   �0@��a�n`�?�             o@T       _                    �?4���C�?            �@@U       ^                    -@����X�?
             ,@V       W                    �?���Q��?             $@������������������������       �                      @X       ]                    @      �?              @Y       \                   P2@և���X�?             @Z       [                    #@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @`       g                    @���y4F�?             3@a       b                    �?և���X�?             @������������������������       �                      @c       d                    �?���Q��?             @������������������������       �                      @e       f                 032@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@i       �                    �?��ݼ��?�            �j@j       {                    �? 1_#�?)            �M@k       n                    �?X�<ݚ�?             2@l       m                    �?      �?              @������������������������       �                     �?������������������������       �                     �?o       z                 pF @     ��?
             0@p       q                    4@X�Cc�?	             ,@������������������������       �                     �?r       s                 �|�9@�	j*D�?             *@������������������������       �                     �?t       y                    �?�q�q�?             (@u       v                 ���@�����H�?             "@������������������������       �                      @w       x                 �&B@؇���X�?             @������������������������       �r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @|       }                 ���@� ��1�?            �D@������������������������       �                     @~       �                    �?������?             A@       �                    �?��a�n`�?             ?@�       �                 ��*@�q�q�?             8@�       �                    �?��+7��?             7@�       �                   @8@      �?              @������������������������       �                     �?�       �                   @@����X�?             @�       �                 �|=@      �?             @������������������������       �                      @������������������������       �      �?              @�       �                    ?@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 �|Y=@z�G�z�?	             .@������������������������       �                     @������������������������       �                     (@������������������������       �                     �?������������������������       �                     @�       �                    >@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?8�Z$���?i            �c@�       �                    �?      �?             B@�       �                    �?�G�z��?             4@�       �                    �?���Q��?             .@�       �                    3@�q�q�?             (@������������������������       �                     @�       �                 pf�@�<ݚ�?             "@�       �                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �|Y>@؇���X�?             @������������������������       �                     @�       �                    A@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 �!@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 X�,@@���Q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        
             0@�       �                    �?      �?P             ^@�       �                 �T)D@��0{9�?@            �W@�       �                 �?�@�)�Db��??            @W@�       �                 �?$@�C��2(�?             F@�       �                   @6@r�q��?             8@������������������������       �                      @�       �                   �8@      �?
             0@������������������������       �                      @�       �                 �|�=@؇���X�?	             ,@�       �                 �|Y=@�q�q�?             @������������������������       �                     @�       �                 ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     4@�       �                 @3�@Jm_!'1�?!            �H@������������������������       �                     @�       �                 pf� @�����H�?            �F@�       �                 ��) @PN��T'�?             ;@�       �                   @F@HP�s��?             9@�       �                    4@ �q�q�?             8@������������������������       �      �?             @������������������������       �                     4@������������������������       �                     �?������������������������       �                      @�       �                 ���"@�X�<ݺ?             2@������������������������       �                     &@�       �                    �?؇���X�?             @�       �                   �<@r�q��?             @������������������������       �                     @�       �                    A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    6@ ��WV�?             :@�       �                    �?�q�q�?             @�       �                 �Y�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@re  trf  bh�h"h#K �rg  h%�rh  Rri  (KK�KK�rj  hR�BP       �q@      d@     �V@     @Z@     �E@     �M@      7@      *@      7@      (@      0@      (@              @      0@       @      .@      @      *@      @      @      @      @      @      @       @      @                       @              @      @              @               @              �?      @              �?      �?       @               @      �?              @                      �?      4@      G@      0@      1@              @      0@      $@       @      $@       @              @      $@              $@      @               @              @      =@      �?      7@              0@      �?      @              @      �?       @      �?                       @      @      @              @      @              H@      G@              "@      H@     �B@      8@      ;@              @      8@      7@              .@      8@       @      .@       @      .@      @      $@      �?      �?      �?              �?      �?              "@              @      @      @               @      @              @       @                       @      "@              8@      $@      8@      "@      @      @      �?      @               @      �?      @      �?                      @      @              4@      @              @      4@                      �?      h@      L@      3@      ,@      @      $@      @      @               @      @      @      @      @      �?      @              @      �?              @                      �?              @      .@      @      @      @               @      @       @       @              �?       @               @      �?              (@             �e@      E@     �D@      2@       @      $@      �?      �?              �?      �?              @      "@      @      "@      �?              @      "@              �?      @       @      �?       @               @      �?      @      �?      @              �?      @               @             �@@       @      @              :@       @      8@      @      1@      @      1@      @      @      @              �?      @       @      @      �?       @              �?      �?       @      �?              �?       @              (@      @              @      (@                      �?      @               @      �?              �?       @             �`@      8@      ;@      "@      &@      "@      "@      @      @      @              @      @       @      �?      �?              �?      �?              @      �?      @              �?      �?              �?      �?               @      �?              �?       @               @      @       @      �?              �?       @                       @      0@             @Z@      .@      T@      ,@      T@      *@      D@      @      4@      @       @              (@      @               @      (@       @      @       @      @              �?       @      �?                       @       @              4@              D@      "@              @      D@      @      7@      @      7@       @      7@      �?      @      �?      4@                      �?               @      1@      �?      &@              @      �?      @      �?      @              �?      �?              �?      �?              �?                      �?      9@      �?       @      �?      �?      �?      �?                      �?      �?              7@        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B8*         4                    �?N9�U-�?           �{@       3                    @��}*_��?1            @T@                           �?      �?0             T@       	                    4@�MI8d�?            �B@                             @      �?              @������������������������       �                     �?                          �0@և���X�?             @������������������������       �                     @������������������������       �                     @
                            @ 	��p�?             =@������������������������       �                     6@                        ���%@����X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       2                    �?�+��<��?            �E@       )                 ���=@��6���?             E@                            �?���Q��?             9@������������������������       �                     �?       &                    �?�q�q�?             8@                            @     ��?             0@                        ���,@      �?              @������������������������       �                     �?������������������������       �                     �?       %                    �?և���X�?	             ,@       $                 xF*@�q�q�?             (@                        ���@z�G�z�?             $@������������������������       �                      @                          �5@      �?              @������������������������       �                     �?        !                 �|�:@؇���X�?             @������������������������       �                      @"       #                 �|�=@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @'       (                     @      �?              @������������������������       �                     �?������������������������       �                     @*       1                 �̾w@������?             1@+       0                     �?     ��?
             0@,       -                 X�lE@���!pc�?             &@������������������������       �                     @.       /                   `P@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?5       `                 `�X!@�ՁE�?�            �v@6       7                 pff@��v����?U            �`@������������������������       �                     8@8       I                    �?�2����?E            �[@9       H                    �?|��?���?             ;@:       A                    9@      �?             :@;       <                 �&B@X�Cc�?             ,@������������������������       �                      @=       @                   �3@r�q��?             @>       ?                   �0@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @B       G                    �?�q�q�?             (@C       F                 `f�@�q�q�?             @D       E                  s�@z�G�z�?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?J       ]                   �E@ ,U,?��?5            �T@K       T                 �?�@H�!b	�?3            @T@L       M                 �|Y<@ pƵHP�?             J@������������������������       �                     :@N       S                 �|�=@ ��WV�?             :@O       P                    �?�IєX�?             1@������������������������       �                     *@Q       R                  sW@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@U       X                 @3�@ܷ��?��?             =@V       W                    �?���Q��?             @������������������������       �                      @������������������������       �                     @Y       \                   �3@ �q�q�?             8@Z       [                    2@r�q��?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     2@^       _                 @3�@      �?              @������������������������       �                     �?������������������������       �                     �?a       |                    �?�zӟ|�?�            �l@b       w                    �?���c��?<            �W@c       l                     @     ��?3             T@d       k                    �? pƵHP�?#             J@e       f                     �? 7���B�?             ;@������������������������       �                     .@g       h                    �?�8��8��?	             (@������������������������       �                     "@i       j                    D@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     9@m       n                 @3�"@      �?             <@������������������������       �                     @o       p                    @�û��|�?             7@������������������������       �                     @q       r                   �:@�d�����?             3@������������������������       �                      @s       v                 ���4@�eP*L��?             &@t       u                 ���$@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @x       {                    @�r����?	             .@y       z                 �̤=@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@}       �                     �?6kh�h��?Z            �`@~       �                   �F@��+��?            �B@       �                   �@@�X����?             6@�       �                    �?և���X�?	             ,@�       �                    �?�eP*L��?             &@�       �                 �|Y>@և���X�?             @�       �                    <@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                 `f�K@      �?             @������������������������       �                      @������������������������       �                      @�       �                 ���i@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �C@      �?              @������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?�       �                  x#J@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   @J@z�G�z�?             .@�       �                    �?      �?              @�       �                 `f�;@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?B�1V���?A            @X@�       �                    �?b:�&���?7            �T@�       �                    &@�r����?'             N@�       �                    5@�q�q�?             (@������������������������       �                     @�       �                     @�����H�?             "@������������������������       �                     @�       �                   �"@z�G�z�?             @������������������������       �                     @�       �                   �<@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    ?@�8��8��?             H@������������������������       �                     9@�       �                     @�㙢�c�?             7@�       �                   @A@@�0�!��?	             1@�       �                    1@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                 `f�)@�8��8��?             (@������������������������       �                     @�       �                   @D@      �?              @������������������������       �                     @�       �                    G@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?r�q��?             @�       �                   �A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     @8����?             7@�       �                    &@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    )@�θ�?             *@������������������������       �                     @������������������������       �                     $@������������������������       �        
             ,@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B       0q@      e@      >@     �I@      >@      I@      @      ?@      @      @              �?      @      @              @      @               @      ;@              6@       @      @              @       @      �?       @                      �?      8@      3@      7@      3@      $@      .@              �?      $@      ,@      "@      @      �?      �?              �?      �?               @      @       @      @       @       @       @              @       @              �?      @      �?       @              @      �?       @      �?       @                       @               @      �?      @      �?                      @      *@      @      *@      @       @      @      @              @      @              @      @              @                      �?      �?                      �?     �n@     �]@      ]@      2@      8@              W@      2@      ,@      *@      *@      *@      @      "@               @      @      �?       @      �?       @                      �?      @               @      @       @      @      �?      @              �?      �?      @      �?              @              �?             �S@      @     @S@      @     �I@      �?      :@              9@      �?      0@      �?      *@              @      �?              �?      @              "@              :@      @      @       @               @      @              7@      �?      @      �?      @              �?      �?      2@              �?      �?              �?      �?              `@      Y@      <@     �P@      .@     @P@      �?     �I@      �?      :@              .@      �?      &@              "@      �?       @               @      �?                      9@      ,@      ,@              @      ,@      "@              @      ,@      @       @              @      @       @      @       @                      @      @              *@       @      @       @      @                       @      $@             @Y@     �@@      3@      2@      @      .@      @       @      @      @      @      @      �?      @      �?                      @       @               @       @       @                       @      �?       @               @      �?              �?      @              @      �?      @              �?      �?      @      �?                      @      (@      @      @      @      @      @              @      @               @              @             �T@      .@      Q@      .@      J@       @       @      @              @       @      �?      @              @      �?      @              �?      �?      �?                      �?      F@      @      9@              3@      @      ,@      @      @       @               @      @              &@      �?      @              @      �?      @               @      �?              �?       @              @      �?      �?      �?              �?      �?              @              0@      @      @      @              @      @              $@      @              @      $@              ,@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B�         t                 ��H@R��O�?           �{@       #                    �??Z���?�            x@                          P,@����?<            @V@                        @�"@��Hg���?            �F@                           �?d��0u��?             >@                          �4@����"�?             =@       
                    �?z�G�z�?             @       	                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                         ��@�q�q�?             8@                           �?�KM�]�?             3@������������������������       �        
             1@������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �        
             .@       "                    @�eP*L��?              F@                            @�n_Y�K�?            �C@������������������������       �                     4@       !                    @���y4F�?             3@                           @�t����?             1@                           �?��S�ۿ?             .@������������������������       �                     @                        ���5@      �?              @                        X�,@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                            @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @$       1                     �?���I�?�            �r@%       0                   @M@�n_Y�K�?             :@&       '                 ��$:@�G��l��?             5@������������������������       �                      @(       /                    H@�θ�?             *@)       .                   �>@�z�G��?             $@*       -                 ��=@      �?              @+       ,                 `f�;@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @2       G                     @��0k��?�            �p@3       F                   �3@8�Z$���?&            @P@4       9                    �?�GN�z�?             F@5       6                 �|Y:@      �?             @������������������������       �                      @7       8                 ���,@      �?              @������������������������       �                     �?������������������������       �                     �?:       E                   �+@R���Q�?             D@;       @                 �|Y=@�MI8d�?            �B@<       ?                    &@�IєX�?             1@=       >                    5@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@A       B                 `f�)@      �?             4@������������������������       �                      @C       D                   �A@�q�q�?             (@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �        
             5@H       [                    �?�M��?y            �i@I       Z                    �?:ɨ��?            �@@J       K                 ���@�������?             >@������������������������       �                     @L       S                 �|Y=@8����?             7@M       R                    �?�eP*L��?             &@N       O                   @@�q�q�?             "@������������������������       �                     @P       Q                   �2@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @T       Y                 �|Y?@r�q��?             (@U       X                    �?�<ݚ�?             "@V       W                   @@�q�q�?             @������������������������       ����Q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @\       s                    �?���@�c�?f            �e@]       ^                    �?������?Z            �b@������������������������       �                     7@_       `                    #@     ��?K             `@������������������������       �                     �?a       d                 `f�@��b�h8�?J            �_@b       c                    6@�q�q�?             @������������������������       �                      @������������������������       �                     �?e       f                 �?�@�&/�E�?H             _@������������������������       �                     I@g       h                 @3�@�����?,            �R@������������������������       �                     @i       r                    �?����Q8�?*            �Q@j       k                   �0@�>����?              K@������������������������       �      �?              @l       q                 pf� @0G���ջ?             J@m       p                 ��) @��a�n`�?             ?@n       o                    4@XB���?             =@������������������������       ��q�q�?             @������������������������       �                     :@������������������������       �                      @������������������������       �                     5@������������������������       �        
             1@������������������������       �                     5@u       x                    �?�e�,��?*            �M@v       w                    @Pa�	�?            �@@������������������������       �                     @@������������������������       �                     �?y       |                 �D�M@�	j*D�?             :@z       {                 0�"K@�q�q�?             @������������������������       �                      @������������������������       �                     @}       �                    �?z�G�z�?             4@~       �                     �?      �?              @       �                    C@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �1@      �?	             (@������������������������       �                     �?�       �                 X�l@@"pc�
�?             &@������������������������       �                     @�       �                   @E@�q�q�?             @������������������������       �                     �?�       �                 03�S@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B�       0s@      a@      r@     @X@      ?@      M@      &@      A@      &@      3@      &@      2@      @      �?       @      �?       @                      �?       @              @      1@       @      1@              1@       @              @                      �?              .@      4@      8@      .@      8@              4@      .@      @      .@       @      ,@      �?      @              @      �?      @      �?      @                      �?      @              �?      �?              �?      �?                       @      @             p@     �C@      0@      $@      &@      $@       @              @      $@      @      @      �?      @      �?      @              @      �?                      @       @                      @      @              n@      =@     �K@      $@      A@      $@      @      �?       @              �?      �?              �?      �?              ?@      "@      ?@      @      0@      �?      @      �?              �?      @              &@              .@      @       @              @      @              @      @                      @      5@             @g@      3@      7@      $@      7@      @      @              0@      @      @      @      @      @      @              @      @      @                      @               @      $@       @      @       @      @       @      @       @      �?              @              @                      @     `d@      "@     �a@      "@      7@             �]@      "@              �?     �]@       @       @      �?       @                      �?     @]@      @      I@             �P@      @              @     �P@      @      I@      @      �?      �?     �H@      @      <@      @      <@      �?       @      �?      :@                       @      5@              1@              5@              3@      D@      �?      @@              @@      �?              2@       @       @      @       @                      @      0@      @      @      �?      @      �?      @                      �?       @              "@      @              �?      "@       @      @              @       @              �?      @      �?      �?      �?      �?                      �?      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B�$                             �?�r*e���?           �{@������������������������       �                     "@       �                  x#J@z�Q�/�?           0{@       }                    �?8�{�?�            �v@       *                    �?
v��?�            �t@                            @�q�Q�?<             X@                         ��9@�?�|�?            �B@������������������������       �                     3@	       
                    �?�X�<ݺ?             2@������������������������       �                     @                           �?��S�ۿ?
             .@                           D@؇���X�?             @������������������������       �                     @                        `ff@@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                        ��@��Q:��?!            �M@������������������������       �        	             2@                           �?D^��#��?            �D@                           �?և���X�?             @                        P��+@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @       )                 �̼6@�ʻ����?             A@       $                    �?X�<ݚ�?             ;@       !                    �?�ՙ/�?             5@                           �?���|���?	             &@������������������������       �                     �?                         `�X!@���Q��?             $@������������������������       �                     @������������������������       �                     @"       #                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?%       &                 �!@�q�q�?             @������������������������       �                     �?'       (                 ��,2@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @+       B                 �?�@�uD����?�             m@,       ;                    �?t��ճC�?=             V@-       .                 ���@�>4և��?             <@������������������������       �                     @/       8                 03s@��<b���?             7@0       7                 ��(@z�G�z�?             4@1       6                 �|Y=@���y4F�?             3@2       5                    �?�q�q�?             @3       4                   �5@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@������������������������       �                     �?9       :                 �|Y=@�q�q�?             @������������������������       �                     �?������������������������       �                      @<       A                    @ �.�?Ƞ?%             N@=       >                     @�8��8��?             (@������������������������       �                      @?       @                    6@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     H@C       D                    !@ ]�к��?^             b@������������������������       �                      @E       F                 @3�@"pc�
�?\            �a@������������������������       �                     @G       V                     �?*
;&���?Y            @a@H       U                   @M@��Q��?             4@I       T                 0�E@j���� �?             1@J       K                 ��$:@���|���?	             &@������������������������       �                     �?L       O                    �?�z�G��?             $@M       N                 X�lE@      �?              @������������������������       �                     �?������������������������       �                     �?P       Q                 `f�;@      �?              @������������������������       �                     @R       S                 X��B@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @W       |                 �y�/@�^����?I            �]@X       w                    �?�T|n�q�?6            �U@Y       v                   �+@��r�Z}�?3            �S@Z       ]                   �0@b�h�d.�?.            �Q@[       \                    �?      �?             @������������������������       ��q�q�?             @������������������������       �                     �?^       k                 �|Y=@��2(&�?+            �P@_       d                 ���$@�˹�m��?             C@`       c                   �3@`2U0*��?             9@a       b                 pf� @r�q��?             @������������������������       �      �?              @������������������������       �                     @������������������������       �        	             3@e       j                    4@8�Z$���?
             *@f       g                   �2@���Q��?             @������������������������       �                      @h       i                   �'@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @l       o                 �|>@d}h���?             <@m       n                 ��) @      �?             $@������������������������       �                     @������������������������       �                     @p       u                 pf� @�X�<ݺ?             2@q       r                   @F@؇���X�?             @������������������������       �                     @s       t                    I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             &@������������������������       �                     "@x       y                    �?����X�?             @������������������������       �                     �?z       {                 �=/@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @@~                            @�C��2(�?            �@@������������������������       �                     @������������������������       �                     >@�       �                 �|�=@�Jhu4��?(            @R@�       �                    :@�q�q�?             >@�       �                    �?��.k���?             1@�       �                    �?X�Cc�?             ,@������������������������       �                     @�       �                    �?X�<ݚ�?             "@�       �                   �5@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �4@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                 p�O@8�Z$���?             *@������������������������       �                     �?�       �                    �?�8��8��?             (@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                 03�S@>��C��?            �E@�       �                 03�M@���}<S�?             7@������������������������       �                     "@�       �                    �?؇���X�?	             ,@������������������������       �                     "@�       �                    �?���Q��?             @�       �                 8�<Q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?���Q��?             4@������������������������       �                     @�       �                    �?��S���?             .@������������������������       �                     @�       �                    �?�q�q�?             (@������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�Bp
       �q@     @d@              "@     �q@      c@     �o@     �[@     �k@     �Z@      7@     @R@      �?      B@              3@      �?      1@              @      �?      ,@      �?      @              @      �?       @      �?                       @               @      6@     �B@              2@      6@      3@      @      @      @       @               @      @                       @      3@      .@      (@      .@       @      *@      @      @      �?              @      @      @                      @      �?      "@              "@      �?              @       @              �?      @      �?      @                      �?      @             �h@      A@     �T@      @      7@      @      @              2@      @      0@      @      .@      @       @      @       @      �?              �?       @                      @      *@              �?               @      �?              �?       @             �M@      �?      &@      �?       @              @      �?      @                      �?      H@             @]@      <@               @     @]@      :@              @     @]@      5@      *@      @      $@      @      @      @      �?              @      @      �?      �?      �?                      �?       @      @              @       @      @              @       @              @              @              Z@      ,@      R@      ,@     �P@      (@      M@      (@      �?      @      �?       @              �?     �L@      "@     �A@      @      8@      �?      @      �?      �?      �?      @              3@              &@       @      @       @       @              �?       @               @      �?               @              6@      @      @      @      @                      @      1@      �?      @      �?      @              �?      �?              �?      �?              &@              "@              @       @      �?              @       @      @                       @      @@              >@      @              @      >@              >@     �E@      4@      $@      "@       @      "@      @      @              @      @       @      @       @                      @       @       @       @                       @              @      &@       @              �?      &@      �?      @      �?              �?      @              @              $@     �@@       @      5@              "@       @      (@              "@       @      @      �?      �?      �?                      �?      �?       @      �?                       @       @      (@              @       @      @              @       @      @              @       @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B8*         $                    �?�K�n���?           �{@       	                    �?և���X�?0            @S@                           �?      �?             @@������������������������       �                     :@                           �?r�q��?             @                             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @
       #                    �?���X�K�?            �F@                           �?�^�����?            �E@                          �8@��R[s�?            �A@������������������������       �                     "@                           �?$��m��?             :@                            �?��H�}�?             9@                          �O@�q�q�?             (@                        X�lC@      �?              @                        ��2>@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                        �|Y=@�	j*D�?             *@������������������������       �                     @������������������������       �                     "@������������������������       �                     �?                        ԼGC@      �?              @������������������������       �                     @                           >@z�G�z�?             @������������������������       �                      @       "                    �?�q�q�?             @        !                 ڪ�q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @%       \                     @�+:���?�            �v@&       A                    �?��`�K�?Y            `c@'       *                    �?`Y���?5            �V@(       )                   �'@ 	��p�?             =@������������������������       �                      @������������������������       �                     ;@+       @                   @J@¦	^_�?#             O@,       ?                   �>@ҳ�wY;�?            �I@-       4                     �?��
ц��?            �C@.       /                   �B@��Q��?             4@������������������������       �                     @0       1                 �̌*@��
ц��?             *@������������������������       �                     @2       3                 `f�;@؇���X�?             @������������������������       �                     @������������������������       �                     �?5       6                    @�d�����?             3@������������������������       �                     @7       8                    &@     ��?             0@������������������������       �                     �?9       >                   @D@������?
             .@:       ;                 �|�<@8�Z$���?	             *@������������������������       �                     @<       =                   �A@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     (@������������������������       �                     &@B       K                    �?     ��?$             P@C       J                   �:@      �?             @@D       I                     @      �?              @E       H                    �?����X�?             @F       G                    A@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@L       O                   �3@     ��?             @@M       N                    *@����X�?             @������������������������       �                      @������������������������       �                     @P       U                  x�F@��H�}�?             9@Q       R                    �?r�q��?             (@������������������������       �                     @S       T                    :@�q�q�?             @������������������������       �                      @������������������������       �                     @V       W                  x�O@��
ц��?             *@������������������������       �                     @X       [                     �?���Q��?             $@Y       Z                   �I@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @]       �                 �|�=@�T`�[k�?�            �j@^       �                    �?���!pc�?h            �d@_       �                    �?�8�G�V�?W             a@`       �                 �!&B@��i#[�?O            �_@a       h                   �0@������?M            �^@b       c                    �?����X�?             @������������������������       �                     �?d       e                 pf�@�q�q�?             @������������������������       �                     �?f       g                    �?z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @i       x                   �4@&d���?H             ]@j       k                    �?���|���?             6@������������������������       �                      @l       s                   �3@�z�G��?             4@m       n                   �2@؇���X�?             ,@������������������������       �                     @o       p                 �?�@z�G�z�?             $@������������������������       �                     @q       r                 `�8"@�q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @t       u                 @3�@�q�q�?             @������������������������       �                     �?v       w                 pf&!@z�G�z�?             @������������������������       �                     @������������������������       �                     �?y       �                    �?@�҇��?;            �W@z       {                   �7@�P�*�?             ?@������������������������       �                     @|       }                    ;@X�Cc�?             <@������������������������       �                      @~       �                 `�j@�n_Y�K�?             :@       �                 �|Y=@�q�q�?             8@������������������������       �                     �?�       �                 ���@8����?             7@������������������������       �                     @�       �                 ��(@��Q��?             4@�       �                 ���@b�2�tk�?             2@�       �                 ��@      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?X�Cc�?	             ,@������������������������       �r�q��?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?��d��?(            �O@�       �                    �?      �?              @�       �                 pf�@����X�?             @�       �                 pf�@�q�q�?             @������������������������       �                     �?�       �                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?t�6Z���?!            �K@�       �                 �&B@ZՏ�m|�?            �H@�       �                   �@j���� �?             1@������������������������       �                     �?�       �                    7@      �?             0@������������������������       �                     @�       �                   �:@���Q��?             $@������������������������       �                     @�       �                 ��@և���X�?             @������������������������       �                      @�       �                 �|Y=@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                 ���"@      �?             @@������������������������       �                     4@�       �                 ���(@�8��8��?             (@�       �                   �<@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                 032@���Q��?             $@�       �                 �|Y<@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     =@�       �                    �?=QcG��?             �G@�       �                    �?؇���X�?             @������������������������       �                     @�       �                 ���@@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 @3�@P���Q�?             D@�       �                   �C@�r����?
             .@�       �                    C@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     9@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B       pp@     �f@     �@@      F@      �?      ?@              :@      �?      @      �?      �?              �?      �?                      @      @@      *@      >@      *@      :@      "@      "@              1@      "@      0@      "@      @      @      @      @      @      �?              �?      @                      @      @              "@      @              @      "@              �?              @      @              @      @      �?       @               @      �?      �?      �?      �?                      �?      �?               @             �l@      a@     �P@     @V@      G@     �F@       @      ;@       @                      ;@      F@      2@     �@@      2@      5@      2@      @      *@              @      @      @      @              �?      @              @      �?              ,@      @      @              &@      @              �?      &@      @      &@       @      @              @       @               @      @                       @      (@              &@              4@      F@       @      >@       @      @       @      @       @      �?              �?       @                      @              �?              8@      2@      ,@       @      @       @                      @      0@      "@      $@       @      @              @       @               @      @              @      @              @      @      @      @      @              @      @               @             �d@      H@      ^@     �F@     �V@     �F@     �U@     �C@     �U@      B@       @      @              �?       @      @      �?              �?      @               @      �?       @     @U@      ?@      ,@       @               @      ,@      @      (@       @      @               @       @      @              @       @      �?       @      @               @      @      �?              �?      @              @      �?             �Q@      7@      2@      *@              @      2@      $@       @              0@      $@      0@       @              �?      0@      @      @              *@      @      &@      @       @       @       @      �?              �?       @                      �?      "@      @      �?      @       @               @                       @     �J@      $@      @       @      @       @      �?       @              �?      �?      �?              �?      �?              @              �?             �G@       @     �D@       @      $@      @              �?      $@      @      @              @      @              @      @      @       @               @      @       @                      @      ?@      �?      4@              &@      �?      @      �?      @                      �?      @              @                      @      @      @      �?      @              @      �?              @              =@              F@      @      @      �?      @              �?      �?              �?      �?              C@       @      *@       @      @       @      @                       @      @              9@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r   (hKhfK�hgh"h#K �r  h%�r  Rr  (KK��r  hn�B('                             @�/e�U��?           �{@                           @d��0u��?             >@������������������������       �                     1@                           �?8�Z$���?             *@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@	       :                    �?~j`�z�?           �y@
       '                    �?Υf���?)            �N@                           �?��J�fj�?            �B@                          �4@ףp=
�?             $@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                        �|Y=@������?             ;@                        �!�E@      �?             @������������������������       �                     @������������������������       �                     @                             @��s����?             5@                          �O@�z�G��?             $@                            �?      �?             @                        p�w@���Q��?             @                           �?      �?             @                        X�lE@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @!       "                 ���@�C��2(�?             &@������������������������       �                     @#       &                 �|Y?@r�q��?             @$       %                   @@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @(       -                   �7@      �?             8@)       ,                    �?؇���X�?             @*       +                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @.       3                    �?��.k���?             1@/       2                 �|Y>@      �?              @0       1                     @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @4       9                   @K@�<ݚ�?             "@5       8                     �?      �?              @6       7                 ��3Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?;       �                    �?�A kP�?�            v@<       _                    �?p]��t�?�            Pt@=       ^                    @̠�4��?2            �T@>       ]                 0#
9@��Sݭg�?0            �S@?       D                    �?���Q��?             I@@       A                 `f�@�����H�?             "@������������������������       �                     @B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?E       R                 ���&@D^��#��?            �D@F       G                 ���@�����?             3@������������������������       �                     @H       K                 �&B@     ��?             0@I       J                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?L       Q                    �?؇���X�?
             ,@M       N                 `�X!@r�q��?             (@������������������������       �                      @O       P                   �F@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @S       X                    �?���!pc�?
             6@T       U                    �?�θ�?             *@������������������������       �                      @V       W                 03[1@���Q��?             @������������������������       �                      @������������������������       �                     @Y       Z                    �?�q�q�?             "@������������������������       �                     @[       \                     @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@������������������������       �                     @`       �                    �?�y)|���?�            @n@a       b                   �0@��4k��?u            �g@������������������������       �                      @c       �                    �?��C�/��?t            `g@d       �                 ��$:@0��,�?q            �f@e       �                   �D@�J��_��?c            �c@f       m                   �7@��X�-�?W            `a@g       h                 �?�@`Ql�R�?            �G@������������������������       �                     <@i       j                   �2@�}�+r��?
             3@������������������������       �                      @k       l                 pf� @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@n       w                     @���}<S�?@             W@o       p                     �? �q�q�?             8@������������������������       �                     @q       r                 �|Y>@�X�<ݺ?             2@������������������������       �                      @s       v                    @@ףp=
�?             $@t       u                   �'@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @x       y                    �?ДX��?/             Q@������������������������       �                     6@z       �                 �|Y=@*
;&���?!             G@{       �                   �<@������?             1@|                          �8@8�Z$���?	             *@}       ~                   �@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `!@      �?             @������������������������       �                      @������������������������       �                      @�       �                  sW@ܷ��?��?             =@�       �                 pf�@      �?             @������������������������       �                      @������������������������       �                      @�       �                 @3�@`2U0*��?             9@�       �                    B@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�       �                    G@      �?             4@�       �                   @E@      �?             $@������������������������       �                     �?�       �                 ���@X�<ݚ�?             "@������������������������       �                     @�       �                 @3�@�q�q�?             @������������������������       �                     @�       �                   @F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�       �                     @\X��t�?             7@�       �                   �I@�G��l��?             5@�       �                     �?������?	             .@�       �                 `f�;@d}h���?             ,@������������������������       �                     $@�       �                 X��B@      �?             @�       �                   �>@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                     �?�&=�w��?!            �J@�       �                    �?8�Z$���?             *@�       �                   @B@ףp=
�?             $@�       �                 `f�K@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     D@�       �                 ���Y@h�����?             <@������������������������       �                     ;@������������������������       �                     �?r  tr  bh�h"h#K �r  h%�r  Rr	  (KK�KK�r
  hR�B0        s@     �a@      &@      3@              1@      &@       @      �?       @      �?                       @      $@             Pr@     @^@      >@      ?@      5@      0@      �?      "@      �?      �?              �?      �?                       @      4@      @      @      @              @      @              1@      @      @      @      @      @      @       @      @      �?       @      �?       @                      �?      �?                      �?              �?      @              $@      �?      @              @      �?      @      �?       @      �?      �?               @              "@      .@      �?      @      �?      @              @      �?                      @       @      "@      �?      @      �?      @              @      �?                      @      @       @      @      �?       @      �?              �?       @              @                      �?     pp@     �V@     �m@     @V@      9@      M@      4@      M@      4@      >@      �?       @              @      �?      �?      �?                      �?      3@      6@      *@      @              @      *@      @      �?      �?              �?      �?              (@       @      $@       @       @               @       @               @       @               @              @      0@      @      $@               @      @       @               @      @              @      @              @      @      �?              �?      @                      <@      @             `j@      ?@      d@      =@               @      d@      ;@     `c@      ;@      b@      ,@     @`@      "@      G@      �?      <@              2@      �?       @              $@      �?              �?      $@              U@       @      7@      �?      @              1@      �?       @              "@      �?      �?      �?      �?                      �?       @             �N@      @      6@             �C@      @      *@      @      &@       @      @       @               @      @              @               @       @       @                       @      :@      @       @       @       @                       @      8@      �?      @      �?      @                      �?      2@              .@      @      @      @              �?      @      @      @               @      @              @       @      �?       @                      �?      $@              $@      *@      $@      &@      @      &@      @      &@              $@      @      �?      �?      �?              �?      �?               @              �?              @                       @      @             �I@       @      &@       @      "@      �?      @      �?      @                      �?      @               @      �?              �?       @              D@              ;@      �?      ;@                      �?r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfK�hgh"h#K �r!  h%�r"  Rr#  (KKۅr$  hn�B�/         X                    �?��_����?            �{@       W                    @�|�ʒ�?e             c@       H                 Ь�9@z�c�@-�?b            �b@       ?                   @B@h�n��?8            @U@                            @�M;q��?2            �R@������������������������       �                     *@                            �?f���M�?*             O@                        pF @������?             >@	       
                 03�@�㙢�c�?             7@������������������������       �                     �?                        �|�9@��2(&�?             6@������������������������       �                     @                           �?r�q��?
             2@                           �?�t����?	             1@������������������������       �                     @                        ���@r�q��?             (@������������������������       �                      @                        �&B@z�G�z�?             $@������������������������       ��<ݚ�?             "@������������������������       �                     �?������������������������       �                     �?                           �?և���X�?             @                        83�0@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        �|�>@      �?             @                           �?�q�q�?             @                        P�h2@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?!       6                 �|Y<@     ��?             @@"       3                    �?�q�q�?             8@#       .                    �?�����?             3@$       %                 ���@X�<ݚ�?             "@������������������������       �                      @&       '                    3@����X�?             @������������������������       �                     �?(       )                    5@r�q��?             @������������������������       �                      @*       -                 جJ"@      �?             @+       ,                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @/       0                    �?ףp=
�?             $@������������������������       �                     @1       2                 (C�1@�q�q�?             @������������������������       �                      @������������������������       �                     �?4       5                 ��;+@���Q��?             @������������������������       �                     @������������������������       �                      @7       >                     @      �?              @8       =                    �?�q�q�?             @9       <                    �?      �?             @:       ;                 ��� @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @@       E                    �?�z�G��?             $@A       B                   �E@      �?              @������������������������       �                     @C       D                    (@      �?             @������������������������       �                      @������������������������       �                      @F       G                 ��<0@      �?              @������������������������       �                     �?������������������������       �                     �?I       P                    �?$Q�q�?*            �O@J       K                   �E@��<b�ƥ?             G@������������������������       �                     A@L       M                    �?�8��8��?	             (@������������������������       �                     @N       O                   @F@؇���X�?             @������������������������       �                     �?������������������������       �                     @Q       R                    �?@�0�!��?             1@������������������������       �                     @S       T                     @d}h���?	             ,@������������������������       �                     $@U       V                 ��p@@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @Y       x                    �?�&����?�            @r@Z       w                    �?      �?             D@[       p                    �?�d�����?             C@\       i                 ���:@�'�`d�?            �@@]       h                    �?�t����?             1@^       _                 �|=@      �?
             0@������������������������       �                     @`       g                 �|�=@z�G�z�?             $@a       b                     @����X�?             @������������������������       �                     �?c       d                 ���@�q�q�?             @������������������������       �                     �?e       f                   @@���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?j       k                 @�@@     ��?             0@������������������������       �                     @l       m                 ��hU@8�Z$���?             *@������������������������       �                     @n       o                 p"�X@�q�q�?             @������������������������       �                      @������������������������       �                     @q       t                    �?���Q��?             @r       s                ��k(@      �?              @������������������������       �                     �?������������������������       �                     �?u       v                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @y       �                 ���X@0,Tg��?�            �o@z       �                    �?���O1��?�             o@{       �                 �|Y=@HP�s��?             9@|                           �?�<ݚ�?             "@}       ~                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     0@�       �                     �?>4և�z�?�             l@�       �                    �?�z�G��?             D@�       �                    J@�q�q�?             B@�       �                   �G@X�<ݚ�?             ;@�       �                   �F@���Q��?             9@�       �                   �D@�G��l��?             5@�       �                 ��$:@D�n�3�?             3@������������������������       �                     @�       �                    �?�q�q�?	             (@�       �                 �|Y>@      �?              @������������������������       �                     @�       �                   �@@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    9@      �?             @������������������������       �                     �?�       �                   @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                     @�       �                 �G�?�A����?v             g@������������������������       �                     �?�       �                 �?�@Xny��?u            �f@�       �                     @P����?%            �M@������������������������       �                     @�       �                    �?�h����?#             L@�       �                 @3�@���J��?             �I@�       �                    6@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �G@������������������������       �                     @�       �                     @�חF�P�?P             _@�       �                    �?�MI8d�?            �B@�       �                    1@@�0�!��?             A@�       �                   �@@���!pc�?             6@�       �                 `f�&@؇���X�?
             ,@�       �                    5@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                 `fF)@�����H�?             "@������������������������       �                     �?�       �                   �=@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �A@      �?              @������������������������       �                     @�       �                   @D@z�G�z�?             @������������������������       �                     @�       �                   �'@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     @�       �                   �E@��{H�?5            �U@�       �                    �?؇���X�?3             U@�       �                 @3�@     ��?)             P@������������������������       �                     @�       �                    )@f>�cQ�?'            �N@������������������������       �                     @�       �                   �0@x�}b~|�?%            �L@�       �                 ��L,@�q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @�       �                    �?�IєX�?!            �I@�       �                 �|>@t��ճC�?             F@�       �                 �!&B@��a�n`�?             ?@�       �                 ���#@��S�ۿ?             >@�       �                 ���"@���}<S�?             7@�       �                 pf� @P���Q�?             4@�       �                    4@$�q-�?	             *@������������������������       �      �?              @������������������������       �                     &@������������������������       �                     @�       �                   �<@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     @������������������������       �        
             4@�       �                 @3�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KK�KK�r*  hR�B�       �q@     �d@     �B@     �\@     �@@     �\@      =@      L@      6@     �J@              *@      6@      D@       @      6@      @      3@      �?              @      3@              @      @      .@       @      .@              @       @      $@               @       @       @       @      @              �?      �?              @      @       @      �?       @                      �?       @       @      �?       @      �?      �?      �?                      �?              �?      �?              ,@      2@       @      0@      @      *@      @      @               @      @       @              �?      @      �?       @              @      �?      �?      �?              �?      �?               @              �?      "@              @      �?       @               @      �?               @      @              @       @              @       @      @       @       @       @       @      �?       @                      �?              �?       @               @              @      @      @       @      @               @       @       @                       @      �?      �?      �?                      �?      @     �M@      �?     �F@              A@      �?      &@              @      �?      @      �?                      @      @      ,@              @      @      &@              $@      @      �?              �?      @              @             `n@     �H@      >@      $@      <@      $@      :@      @      .@       @      ,@       @      @               @       @      @       @      �?              @       @      �?              @       @       @       @      �?              @              �?              &@      @              @      &@       @      @              @       @               @      @               @      @      �?      �?              �?      �?              �?       @               @      �?               @             �j@     �C@     �j@      B@      7@       @      @       @      �?       @      �?                       @      @              0@             �g@      A@      <@      (@      8@      (@      .@      (@      .@      $@      &@      $@      &@       @      @              @       @       @      @              @       @      @       @                      @       @       @      �?              �?       @      �?                       @               @      @                       @      "@              @             @d@      6@              �?     @d@      5@      M@      �?      @             �K@      �?      I@      �?      @      �?      @                      �?     �G@              @              Z@      4@      ?@      @      <@      @      0@      @      (@       @      @      �?              �?      @               @      �?      �?              @      �?      @                      �?      @      @              @      @      �?      @              �?      �?      �?                      �?      (@              @             @R@      ,@      R@      (@      J@      (@              @      J@      "@              @      J@      @      @       @      �?       @      @              H@      @     �D@      @      <@      @      <@       @      5@       @      3@      �?      (@      �?      �?      �?      &@              @               @      �?       @                      �?      @                      �?      *@              @              4@              �?       @               @      �?                      @r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfK�hgh"h#K �rA  h%�rB  RrC  (KKͅrD  hn�B�,                             @�r*e���?           �{@                           @�S����?             3@������������������������       �                     .@                           @      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @	       H                     �?n?U���?           �z@
       G                   @N@�q�q��?@             X@       B                    �?�X���?<             V@                        0#�9@���|���?6            @S@������������������������       �                     @                          @>@�Y�R_�?2            �Q@                           �?�8��8��?             (@������������������������       �                     @                           �?      �?              @������������������������       �                     �?                        X�l@@؇���X�?             @������������������������       �                     �?������������������������       �                     @       !                  x#J@:���W�?*            �M@                           �?����X�?	             ,@                           �?      �?             @                         ��@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �|Y>@ףp=
�?             $@                          �>@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @"       A                 ���m@��Hg���?!            �F@#       8                    �?�GN�z�?              F@$       1                 ��UT@     ��?             @@%       .                 ���S@���y4F�?             3@&       '                    �?      �?             0@������������������������       �                     (@(       )                 `�iJ@      �?             @������������������������       �                     �?*       +                    9@�q�q�?             @������������������������       �                     �?,       -                   @C@      �?              @������������������������       �                     �?������������������������       �                     �?/       0                 �|�:@�q�q�?             @������������������������       �                      @������������������������       �                     �?2       3                 �_@$�q-�?
             *@������������������������       �                      @4       7                    �?z�G�z�?             @5       6                 0w�a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?9       >                    �?�q�q�?             (@:       ;                    �?���Q��?             @������������������������       �                     �?<       =                   @K@      �?             @������������������������       �                      @������������������������       �                      @?       @                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?C       F                    �?"pc�
�?             &@D       E                   �6@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @I       z                    �?��aV�?�            �t@J       q                   @B@X�Cc�?;            �X@K       V                   �5@:���u��?1            @S@L       U                   �3@      �?             4@M       P                 �y�+@�q�q�?
             .@N       O                 03�@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@Q       T                    �?z�G�z�?             @R       S                    "@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @W       p                    @�S����?$            �L@X       i                    �?؇���X�?#             L@Y       Z                 ��@��G���?            �B@������������������������       �                     "@[       \                   �8@      �?             <@������������������������       �                     @]       ^                   �:@�X����?             6@������������������������       �                      @_       `                 �|Y=@      �?             4@������������������������       �                     @a       h                     @�q�q�?
             .@b       c                    �?�n_Y�K�?	             *@������������������������       �                      @d       g                 �̌"@���!pc�?             &@e       f                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @j       k                 �|Y<@�}�+r��?
             3@������������������������       �                     &@l       o                 м�9@      �?              @m       n                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?r       w                    G@���N8�?
             5@s       v                     @r�q��?             2@t       u                   �3@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@x       y                   �B@�q�q�?             @������������������������       �                     �?������������������������       �                      @{       �                    �?� p�	��?�            �l@|       �                    �?������?             >@}       �                   @@���B���?             :@~                        ���@�C��2(�?             &@������������������������       �                      @�       �                   �5@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                     @������?             .@�       �                 `��,@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                 м;4@�z�G��?             $@�       �                   �:@      �?              @������������������������       �                      @�       �                    �?r�q��?             @�       �                 �|Y=@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                     @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�7A��?~             i@�       �                    �?Ե��,��?e            �d@�       �                  ��@HP�s��?             9@������������������������       �                      @�       �                 �|Y=@�t����?             1@������������������������       �                      @������������������������       �        
             .@�       �                   �0@��27
��?U            `a@������������������������       �      �?             @�       �                   �7@�\�)G�?S            �`@������������������������       �                    �E@�       �                 0��D@��A��?8             W@�       �                     @,sI�v�?6            �V@�       �                    @@��S�ۿ?             >@�       �                 �|�<@�r����?             .@������������������������       �                     @�       �                 �|Y>@�<ݚ�?             "@�       �                    @r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �'@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     .@�       �                   @C@R���Q�?$             N@�       �                   �9@�����H�?            �F@�       �                   �8@�q�q�?             @�       �                   �@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 @33@      �?             @������������������������       �                     �?������������������������       �                     @�       �                 �|�=@$�q-�?            �C@�       �                 ��) @H%u��?             9@�       �                 �?$@���N8�?             5@�       �                 pf�@z�G�z�?             @������������������������       �                     @�       �                 �|Y=@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             0@�       �                 �̜!@      �?             @������������������������       �                     �?�       �                   �<@�q�q�?             @������������������������       �                     �?�       �                 ���(@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@�       �                   �H@������?             .@�       �                 pf&@      �?              @������������������������       �                      @�       �                 ��	0@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                    �B@rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KK�KK�rJ  hR�B�       �q@     @d@      @      0@              .@      @      �?      �?      �?              �?      �?               @             pq@     @b@      C@      M@      >@      M@      <@     �H@      @              6@     �H@      �?      &@              @      �?      @              �?      �?      @      �?                      @      5@      C@      $@      @      �?      @      �?      �?      �?                      �?               @      "@      �?      @      �?              �?      @              @              &@      A@      $@      A@      @      ;@      @      .@       @      ,@              (@       @       @              �?       @      �?      �?              �?      �?              �?      �?               @      �?       @                      �?      �?      (@               @      �?      @      �?      @      �?                      @              �?      @      @      @       @      �?               @       @       @                       @       @      @              @       @              �?               @      "@       @      @              @       @                      @       @              n@      V@     �A@     �O@      3@      M@      $@      $@      @      $@      �?      "@      �?                      "@      @      �?      �?      �?              �?      �?              @              @              "@      H@       @      H@      @      >@              "@      @      5@              @      @      .@       @              @      .@              @      @      $@      @       @       @              @       @      @      �?              �?      @                      @               @      �?      2@              &@      �?      @      �?       @               @      �?                      @      �?              0@      @      .@      @       @      @              @       @              *@              �?       @      �?                       @     �i@      9@      6@       @      5@      @      $@      �?       @               @      �?              �?       @              &@      @      @      �?              �?      @              @      @      @      @               @      @      �?      @      �?              �?      @               @               @              �?      @      �?                      @      g@      1@     `b@      1@      7@       @       @              .@       @               @      .@              _@      .@       @       @     �^@      *@     �E@             �S@      *@     �S@      &@      <@       @      *@       @      @              @       @      @      �?      @                      �?       @      �?       @                      �?      .@             �I@      "@      D@      @      @       @      �?      �?              �?      �?              @      �?              �?      @              B@      @      6@      @      4@      �?      @      �?      @              �?      �?      �?                      �?      0@               @       @              �?       @      �?      �?              �?      �?              �?      �?              ,@              &@      @      @      @       @               @      @              @       @              @                       @     �B@        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfK�hgh"h#K �ra  h%�rb  Rrc  (KKׅrd  hn�B/         `                     @�/��p�?           �{@       9                    �?����?{            �i@                           1@�oS��?K            ``@������������������������       �                     @       (                    G@��rf�B�?H            @_@                           �?$1�l���?;            @Y@������������������������       �                     8@       %                    �?��cv�?*            @S@	                        �|�<@���o,��?'            @R@
                           4@ ��WV�?             :@                           &@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             4@                           �?��V�I��?            �G@                        ���,@      �?             @������������������������       �                     �?                         `6@���Q��?             @������������������������       �                      @                        ��2>@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �'@�>$�*��?            �D@������������������������       �                     *@       "                     �?X�Cc�?             <@       !                   �@@�����?
             3@                         �|Y>@�eP*L��?             &@                          �>@      �?             $@                           <@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @#       $                   @A@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @&       '                    @@      �?             @������������������������       �                      @������������������������       �                      @)       *                   �G@�q�q�?             8@������������������������       �                     @+       0                    �?�d�����?             3@,       /                    �?      �?             @-       .                   �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?1       2                    �?�r����?             .@������������������������       �                     @3       8                   �J@r�q��?             (@4       5                   �H@�q�q�?             @������������������������       �                     �?6       7                   @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@:       O                    �?^��4m�?0            �R@;       B                    �?�4F����?            �D@<       =                     �?�nkK�?             7@������������������������       �        	             ,@>       ?                   �7@�����H�?             "@������������������������       �                     @@       A                   @B@z�G�z�?             @������������������������       �                     @������������������������       �                     �?C       N                   �G@�q�q�?             2@D       I                    �?      �?             0@E       H                   �:@z�G�z�?             @F       G                   �5@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @J       M                 03�M@���!pc�?             &@K       L                  x#J@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @P       ]                    @"pc�
�?            �@@Q       V                     �?�r����?             >@R       S                    H@      �?             (@������������������������       �                      @T       U                    L@      �?             @������������������������       �                     @������������������������       �                     �?W       X                   �8@�X�<ݺ?             2@������������������������       �                     &@Y       \                    =@؇���X�?             @Z       [                 ��A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^       _                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @a       �                    �?
]�YC��?�            �m@b       �                 0�H@���BK�?�            �j@c       j                   �0@��eN_:�?�             j@d       i                    @D�n�3�?             3@e       h                 @� @�8��8��?
             (@f       g                 ���@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @k       �                    �?H~��D
�?v            �g@l       �                    �?���7Qv�?r             g@m       r                    �?���|���?             F@n       o                 ���%@؇���X�?             @������������������������       �                     @p       q                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @s       x                    �?�Gi����?            �B@t       w                    �?X�<ݚ�?             "@u       v                    @r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @y       �                    �?��>4և�?             <@z       {                 �&B@�����?
             3@������������������������       �                      @|       }                 `�X!@�eP*L��?             &@������������������������       �                     @~       �                   �:@r�q��?             @       �                    4@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?X�<ݚ�?             "@�       �                   �3@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                 @3�@��l��?Y            �a@������������������������       �                     �?�       �                   �<@�d�g��?X            �a@�       �                    �?      �?%             P@�       �                   �4@`Jj��?$             O@�       �                    �?�LQ�1	�?             7@�       �                    �?ףp=
�?
             4@������������������������       �                     �?�       �                 ��@�}�+r��?	             3@������������������������       �                     "@�       �                   �3@ףp=
�?             $@�       �                    2@z�G�z�?             @������������������������       �                     �?�       �                 �̌&@      �?             @������������������������       �      �?              @������������������������       �                      @������������������������       �                     @�       �                 �Y�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 ��@ ���J��?            �C@�       �                 ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     B@������������������������       �                      @�       �                    �?h�˹�?3             S@�       �                 �|Y=@�Z��L��?/            �Q@�       �                 ��@      �?             @������������������������       �                     �?�       �                   `!@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�qM�R��?+            �P@�       �                 �|�=@d}h���?	             ,@�       �                 ���@���!pc�?             &@������������������������       �                     @�       �                   @@և���X�?             @������������������������       ����Q��?             @������������������������       �                      @������������������������       �                     @�       �                   @C@ �h�7W�?"            �J@�       �                 �|�=@��Y��]�?            �D@�       �                    �?`2U0*��?             9@�       �                 ��) @ �q�q�?             8@������������������������       �                     4@�       �                 pf� @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        	             0@�       �                   �C@r�q��?             (@������������������������       �                     �?�       �                    �?�C��2(�?             &@������������������������       �                      @�       �                 pf�@�����H�?             "@������������������������       �                     @�       �                   �E@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                  S�-@z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                 ���3@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?$�q-�?             :@������������������������       �                     @�       �                 ��T?@���}<S�?             7@������������������������       �        
             ,@�       �                    �?�<ݚ�?             "@�       �                    @      �?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @re  trf  bh�h"h#K �rg  h%�rh  Rri  (KK�KK�rj  hR�Bp       �p@     �e@     �V@     �\@      R@     �M@              @      R@     �J@     �J@      H@              8@     �J@      8@     �I@      6@      9@      �?      @      �?              �?      @              4@              :@      5@      @      @              �?      @       @       @              �?       @               @      �?              7@      2@      *@              $@      2@      @      *@      @      @      @      @      �?      @      �?                      @      @              �?                       @      @      @              @      @               @       @       @                       @      3@      @      @              ,@      @      �?      @      �?       @      �?                       @              �?      *@       @      @              $@       @      �?       @              �?      �?      �?      �?                      �?      "@              3@     �K@      *@      <@      �?      6@              ,@      �?       @              @      �?      @              @      �?              (@      @      (@      @      @      �?      �?      �?      �?                      �?      @               @      @      @      @      @                      @      @                       @      @      ;@      @      :@      @      "@               @      @      �?      @                      �?      �?      1@              &@      �?      @      �?      �?              �?      �?                      @       @      �?              �?       @             �f@     �M@     �c@     �L@     �c@     �J@       @      &@      �?      &@      �?      @              @      �?                       @      @             �b@      E@     �a@      E@      0@      <@      �?      @              @      �?       @      �?                       @      .@      6@      @      @      �?      @      �?                      @      @              &@      1@      @      *@               @      @      @      @              �?      @      �?       @               @      �?                      @      @      @      @       @               @      @                       @     �_@      ,@              �?     �_@      *@      N@      @      M@      @      4@      @      2@       @              �?      2@      �?      "@              "@      �?      @      �?      �?              @      �?      �?      �?       @              @               @      �?       @                      �?      C@      �?       @      �?       @                      �?      B@               @             �P@      "@     �O@       @       @       @              �?       @      �?       @                      �?     �N@      @      &@      @       @      @      @              @      @       @      @       @              @              I@      @      D@      �?      8@      �?      7@      �?      4@              @      �?              �?      @              �?              0@              $@       @              �?      $@      �?       @               @      �?      @               @      �?       @                      �?      @      �?       @               @      �?      �?              �?      �?              �?      �?              @                      @      8@       @      @              5@       @      ,@              @       @       @       @      �?       @               @      �?              �?              @        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B�%         @                    �?X��d�?�?           �{@       7                    �?t�0i��?W            `a@       6                    @���!pc�?L            @^@                           �?�����?I            @]@                        �|Y:@ �q�q�?             8@������������������������       �                     $@       
                 Pv;@@4և���?             ,@       	                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@       !                 03S$@���U��?:            @W@                            �?d��0u��?             >@                           �?����"�?             =@                         s�@X�<ݚ�?             "@������������������������       �                     @                        �|�9@r�q��?             @������������������������       �                     �?                         s�@z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @                        ���@�z�G��?             4@������������������������       �                     @                         SE"@@�0�!��?             1@                        `�X!@      �?             (@                          �7@ףp=
�?             $@                           5@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?"       %                    �?؇���X�?&            �O@#       $                 �|�>@�q�q�?             @������������������������       �                     �?������������������������       �                      @&       +                    �?�?�P�a�?$             N@'       *                 `f�%@ ���J��?            �C@(       )                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     B@,       3                    �?����X�?             5@-       2                    B@"pc�
�?             &@.       1                    1@ףp=
�?             $@/       0                 `f7@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?4       5                     @���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @8       ?                 �|�=@�<ݚ�?             2@9       :                    @      �?
             0@������������������������       �                     $@;       >                    @�q�q�?             @<       =                 ��T?@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @A       �                  x#J@���gc��?�            s@B       Y                    �?4ԡ"���?�            �p@C       V                    �?f���M�?             ?@D       G                   �5@      �?             8@E       F                    '@�q�q�?             @������������������������       �                     �?������������������������       �                      @H       K                     �?��s����?             5@I       J                 X�lE@      �?             @������������������������       �                     @������������������������       �                     �?L       U                    �?@�0�!��?
             1@M       N                 ���@d}h���?             ,@������������������������       �                     @O       P                 �|�:@�q�q�?             "@������������������������       �                      @Q       T                 �|�=@և���X�?             @R       S                   @@      �?             @������������������������       ����Q��?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @W       X                     @����X�?             @������������������������       �                      @������������������������       �                     @Z       u                 ��) @3e��?�            `m@[       h                 ���@�]��?B            �Y@\       ]                     @�C��2(�?             6@������������������������       �                      @^       g                    ;@؇���X�?
             ,@_       f                    �?�q�q�?             @`       a                    @���Q��?             @������������������������       �                     �?b       c                    �?      �?             @������������������������       �                      @d       e                 ���@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @i       p                    �?F|/ߨ�?2            @T@j       o                 ��@`׀�:M�?-            �R@k       n                 �|Y=@ �q�q�?             8@l       m                    ;@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �        
             ,@������������������������       �                     I@q       t                    �?؇���X�?             @r       s                 pff@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @v       {                    @��2(&�?S            �`@w       x                 �Q��?r�q��?             @������������������������       �                      @y       z                    @      �?             @������������������������       �                     @������������������������       �                     �?|       �                    �?|�(��?N            �_@}       ~                 pf� @@�0�!��?.             Q@������������������������       �                      @       �                 ���"@6YE�t�?-            �P@������������������������       �                     ,@�       �                   �<@���B���?%             J@������������������������       �                     0@�       �                    $@�E��ӭ�?             B@������������������������       �                      @�       �                     @������?             A@�       �                     �?r֛w���?             ?@�       �                   `D@���y4F�?             3@�       �                 ��$:@      �?              @������������������������       �                      @�       �                   �@@�q�q�?             @�       �                 0�?D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@�       �                 `f�)@�q�q�?
             (@������������������������       �                     @�       �                   �3@      �?              @�       �                   �A@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    #@ _�@�Y�?              M@�       �                    !@ףp=
�?             $@������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     H@�       �                   �8@��
ц��?            �C@�       �                     �?     ��?             0@�       �                    �?�q�q�?             (@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                 03�S@8����?             7@�       �                   �I@��S�ۿ?             .@������������������������       �                     &@�       �                   �L@      �?             @������������������������       �                     �?������������������������       �                     @�       �                 @�:x@      �?              @������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B�
       �r@     @b@     �G@      W@     �@@      V@      =@      V@      �?      7@              $@      �?      *@      �?      @              @      �?                      "@      <@     @P@      3@      &@      2@      &@      @      @      @              �?      @              �?      �?      @               @      �?       @      ,@      @              @      ,@      @      "@      @      "@      �?      @      �?      @                      �?      @                       @      @              �?              "@      K@       @      �?              �?       @              @     �J@      �?      C@      �?       @               @      �?                      B@      @      .@       @      "@      �?      "@      �?      @              @      �?                      @      �?              @      @              @      @              @              ,@      @      ,@       @      $@              @       @       @       @       @                       @       @                       @     `o@      K@      m@     �@@      4@      &@      2@      @      �?       @      �?                       @      1@      @      @      �?      @                      �?      ,@      @      &@      @      @              @      @       @              @      @      @      @       @      @      �?              �?              @               @      @       @                      @     �j@      6@     �X@      @      4@       @       @              (@       @      @       @      @       @              �?      @      �?       @              �?      �?      �?                      �?      �?               @             �S@       @     @R@      �?      7@      �?      "@      �?      "@                      �?      ,@              I@              @      �?      @      �?      @                      �?      @             �\@      2@      �?      @               @      �?      @              @      �?             @\@      *@      L@      (@               @      L@      $@      ,@              E@      $@      0@              :@      $@               @      :@       @      7@       @      .@      @      @      @       @               @      @       @      �?              �?       @                      @      &@               @      @      @              @      @      @      @              @      @              �?              @             �L@      �?      "@      �?      @               @      �?              �?       @              H@              2@      5@      &@      @      @      @      @                      @      @              @      0@      �?      ,@              &@      �?      @      �?                      @      @       @      @                       @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B�%         F                     @2��;�O�?           �{@                           �?��S���?y            `h@                          �'@pY���D�?/            �S@������������������������       �                     �?                           �?�(�Tw�?.            �S@                           E@@��8��?             H@������������������������       �                     A@       	                     �?@4և���?             ,@������������������������       �                     &@
                          �3@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     >@                           -@������?J             ]@������������������������       �                     @       !                    �?���GYW�?H            �[@                            �?�r����?             >@                            �?�J�4�?             9@                        �̾w@R���Q�?             4@                           �?�X�<ݺ?             2@������������������������       �                     *@                           �?z�G�z�?             @                        p"4W@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @                        �|Y:@z�G�z�?             @������������������������       �                      @                        ���,@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @"       E                    �?�<ݚ�?6            @T@#       2                 ��$:@�ګH9�?0            �Q@$       %                     �?�?�'�@�?             C@������������������������       �                     @&       1                    �?��hJ,�?             A@'       0                   @A@r�q��?             >@(       -                   �(@�GN�z�?             6@)       ,                    5@$�q-�?	             *@*       +                    &@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@.       /                 �|�<@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @3       >                    �?����e��?            �@@4       =                   �>@�q�q�?             ;@5       6                 03k:@     ��?
             0@������������������������       �                     @7       <                   @=@��
ц��?             *@8       ;                   �J@���|���?             &@9       :                 `f�;@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     &@?       @                 `�iJ@�q�q�?             @������������������������       �                     �?A       D                     �?���Q��?             @B       C                    9@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     $@G       r                    �?΁�)�,�?�             o@H       _                    �?(ǯt��?.            �R@I       ^                    A@��Q��?             D@J       K                 ���@V������?            �B@������������������������       �                     "@L       M                    #@��>4և�?             <@������������������������       �                     @N       W                    �?
;&����?             7@O       R                    �?�z�G��?             $@P       Q                 �|�9@r�q��?             @������������������������       �                     �?������������������������       �z�G�z�?             @S       V                    �?      �?             @T       U                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?X       Y                 ��� @�n_Y�K�?             *@������������������������       �                     @Z       ]                   �8@����X�?             @[       \                 �[$@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @`       q                    @h+�v:�?             A@a       p                   �B@     ��?             @@b       c                    @8�A�0��?             6@������������������������       �                     @d       g                    �?      �?	             2@e       f                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @h       i                    ,@�q�q�?             (@������������������������       �                      @j       o                 м�6@�z�G��?             $@k       l                 �|�>@      �?              @������������������������       �                     @m       n                   �1@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@������������������������       �                      @s       �                 �T�I@�J�4�?l            �e@t       �                 �|Y=@�����	�?i            @e@u       �                    0@��!���?5            @W@v       w                    @p�}�ޤ�?*            @R@������������������������       �                     �?x       �                    �?      �?)             R@y       ~                    �?�'݊U�?&            �P@z       {                 �Y�@�z�G��?             $@������������������������       �                     @|       }                    <@���Q��?             @������������������������       �                      @������������������������       �                     @       �                    �?�k�'7��?!            �L@�       �                   �7@fP*L��?             F@������������������������       �                     7@�       �                 �Y�@�q�q�?             5@�       �                   �8@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                 �̌!@@4և���?	             ,@������������������������       �                     &@�       �                   �<@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 ��Y@�θ�?             *@������������������������       �                     @�       �                 pf�'@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     4@�       �                 �|�=@XI�~�?4            @S@�       �                    �?�����H�?             B@�       �                    �?      �?              @�       �                 ���@r�q��?             @������������������������       �                      @�       �                    �?      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?h�����?             <@�       �                    �?�}�+r��?             3@������������������������       �                     @�       �                 ��) @��S�ۿ?             .@������������������������       �        	             (@�       �                 pf6'@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@�       �                   �E@��Y��]�?            �D@������������������������       �                     A@�       �                   �H@؇���X�?             @�       �                 @3�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B�
       q@     `e@     �V@      Z@       @     @S@      �?              �?     @S@      �?     �G@              A@      �?      *@              &@      �?       @               @      �?                      >@     @V@      ;@              @     @V@      6@      :@      @      5@      @      1@      @      1@      �?      *@              @      �?       @      �?              �?       @               @                       @      @      �?       @               @      �?              �?       @              @             �O@      2@     �J@      2@     �@@      @      @              =@      @      9@      @      1@      @      (@      �?      �?      �?              �?      �?              &@              @      @      @                      @       @              @              4@      *@      2@      "@      @      "@              @      @      @      @      @      �?      @              @      �?              @                       @      &@               @      @              �?       @      @      �?      @      �?                      @      �?              $@             �f@     �P@     �A@     �C@      ,@      :@      &@      :@              "@      &@      1@              @      &@      (@      @      @      �?      @              �?      �?      @       @       @      �?       @      �?                       @      �?               @      @      @               @      @       @       @               @       @                      @      @              5@      *@      3@      *@      "@      *@              @      "@      "@      @       @      @                       @      @      @       @              @      @      �?      @              @      �?       @      �?                       @       @              $@               @             `b@      <@     @b@      8@     �R@      3@      K@      3@              �?      K@      2@      K@      *@      @      @      @               @      @       @                      @     �G@      $@     �B@      @      7@              ,@      @      �?      @              @      �?              *@      �?      &@               @      �?       @                      �?      $@      @      @              @      @              @      @                      @      4@              R@      @      @@      @      @      @      @      �?       @              @      �?       @      �?      �?                       @      ;@      �?      2@      �?      @              ,@      �?      (@               @      �?              �?       @              "@              D@      �?      A@              @      �?      �?      �?              �?      �?              @              �?      @              @      �?        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KKÅr�  hn�B�*         J                     @ �a�e��?           �{@       /                     �?�c:��?s             g@                         x#J@�ɭ�BR�?=            �Y@                        0#�9@��Q���?             D@������������������������       �                     $@                           J@d��0u��?             >@                          `G@D�n�3�?             3@                         �>@և���X�?
             ,@	       
                    �?      �?              @������������������������       �                      @                        ��$:@      �?             @������������������������       �                     �?                        `f�;@���Q��?             @������������������������       �                      @                        X��B@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        �|�9@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@       &                   @I@���N8�?%            �O@                           �?D>�Q�?             J@������������������������       �                     ;@                        03�M@��H�}�?             9@������������������������       �                      @                           �?��.k���?             1@                        �̾w@r�q��?             @������������������������       �                     @������������������������       �                     �?        %                 ��hU@���|���?             &@!       $                    �?z�G�z�?             @"       #                 ���S@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @'       *                    �?�eP*L��?	             &@(       )                 8�tQ@      �?             @������������������������       �                     �?������������������������       �                     @+       .                 `fj@����X�?             @,       -                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @0       9                    �?,ZYN(��?6            @T@1       2                    �?��S�ۿ?             >@������������������������       �                     �?3       8                   @J@ 	��p�?             =@4       5                    E@h�����?             <@������������������������       �                     7@6       7                   @F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?:       I                   �3@�:�]��?!            �I@;       H                    �?\-��p�?             =@<       G                    �?�>����?             ;@=       @                    �?HP�s��?             9@>       ?                 `��,@      �?             @������������������������       �                     �?������������������������       �                     @A       B                 �|Y=@���N8�?             5@������������������������       �                     &@C       D                 `f�)@ףp=
�?	             $@������������������������       �                     @E       F                 X�l@@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �        
             6@K       ~                    �?D'x���?�            @p@L       U                    1@�s��:��?-             S@M       R                    �?      �?	             0@N       O                    �?؇���X�?             @������������������������       �                     @P       Q                    #@      �?              @������������������������       �                     �?������������������������       �                     �?S       T                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?V       ]                    �?�q�q�?$             N@W       X                    5@      �?              @������������������������       �                      @Y       \                 ���0@r�q��?             @Z       [                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^       }                     @���3�E�?             J@_       |                 ���4@�I� �?             G@`       u                    �?\�Uo��?             C@a       r                    �?��X��?             <@b       c                   �4@�	j*D�?             :@������������������������       �                     @d       g                    �?���Q��?             4@e       f                 �&B@      �?             @������������������������       ����Q��?             @������������������������       �                     �?h       k                    8@X�Cc�?             ,@i       j                 جJ"@z�G�z�?             @������������������������       �                     @������������������������       �                     �?l       m                 �|Y>@�����H�?             "@������������������������       �                     @n       o                 ��� @�q�q�?             @������������������������       �                     �?p       q                    A@      �?              @������������������������       �                     �?������������������������       �                     �?s       t                 �|Y<@      �?              @������������������������       �                     �?������������������������       �                     �?v       w                    �?���Q��?             $@������������������������       �                     @x       y                 xFT!@և���X�?             @������������������������       �                      @z       {                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       �                 �T�I@��W���?t             g@�       �                    @�=C|F�?o            �e@�       �                     @��
ц��?	             *@������������������������       �                     @������������������������       �                     @�       �                    �?������?f             d@�       �                 �|Y=@�z�G��?             4@�       �                 �&�)@և���X�?             @������������������������       �                     @�       �                    /@      �?             @������������������������       �                      @�       �                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?8�Z$���?             *@������������������������       �                     &@������������������������       �                      @�       �                 �|Y=@=QcG��?Y            �a@�       �                    �?Xny��?*            �N@�       �                    �?H�ՠ&��?&             K@�       �                    )@L紂P�?#            �I@������������������������       �                     �?�       �                    �?H%u��?"             I@�       �                    �?؇���X�?             E@������������������������       �                     @�       �                 �Y�@�S����?             C@�       �                 @33@�q�q�?             @������������������������       �                     �?�       �                    6@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �3@(N:!���?            �A@�       �                 pf�@      �?	             (@������������������������       �                     @�       �                    2@      �?             @�       �                   �0@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       ��q�q�?             @�       �                   �<@�nkK�?             7@������������������������       �                     5@�       �                 hfF!@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?�(\����?/             T@������������������������       �        
             0@�       �                    �?      �?%             P@�       �                 �?�@@9G��?            �H@������������������������       �                     8@�       �                    �?HP�s��?             9@�       �                   �E@�C��2(�?             6@�       �                 ��) @�X�<ݺ?             2@������������������������       �                     &@�       �                 pf� @؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   �F@      �?             @�       �                 @3�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        	             .@�       �                 p�O@�z�G��?             $@������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�B0        r@     @c@     @W@     �V@      F@     �M@      =@      &@      $@              3@      &@       @      &@       @      @      @      @               @      @      @      �?               @      @               @       @      �?              �?       @              @      �?              �?      @                      @      &@              .@      H@      "@     �E@              ;@      "@      0@               @      "@       @      @      �?      @                      �?      @      @      @      �?       @      �?              �?       @               @                      @      @      @      �?      @      �?                      @      @       @      @       @               @      @               @             �H@      @@       @      <@              �?       @      ;@      �?      ;@              7@      �?      @      �?                      @      �?             �G@      @      9@      @      9@       @      7@       @      @      �?              �?      @              4@      �?      &@              "@      �?      @              @      �?              �?      @               @                       @      6@             �h@     �O@      E@      A@       @      ,@      �?      @              @      �?      �?              �?      �?              �?       @               @      �?              D@      4@      @      @       @              �?      @      �?      �?              �?      �?                      @     �B@      .@      ?@      .@      7@      .@      3@      "@      2@       @      @              (@       @      @      @      @       @              �?      "@      @      �?      @              @      �?               @      �?      @               @      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?              @      @              @      @      @               @      @      �?      @                      �?       @              @             `c@      =@      c@      6@      @      @              @      @             @b@      .@      ,@      @      @      @              @      @      �?       @              �?      �?              �?      �?              &@       @      &@                       @     �`@      "@      K@      @     �G@      @      F@      @              �?      F@      @      B@      @      @              @@      @      �?       @              �?      �?      �?      �?                      �?      ?@      @      "@      @      @              @      @       @      �?      �?      �?      �?              �?       @      6@      �?      5@              �?      �?      �?                      �?       @              @              @             �S@       @      0@              O@       @     �G@       @      8@              7@       @      4@       @      1@      �?      &@              @      �?              �?      @              @      �?      �?      �?              �?      �?               @              @              .@              @      @              @      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfK�hgh"h#K �r�  h%�r�  Rr�  (KK��r�  hn�B�$         (                    �?���&�A�?           �{@       	                    �?���L��?1            �S@                        ���0@ףp=
�?             >@                           �?�z�G��?             $@                           �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     4@
                           �?�q�q�?             H@                        �̾w@�4�����?             ?@                           5@�c�Α�?             =@������������������������       �                     @                        �|Y=@�J�4�?             9@                            @�z�G��?             $@������������������������       �                     @                          @@      �?             @������������������������       �                     @������������������������       �                     @                        X�@@��S�ۿ?	             .@                        4C�2@؇���X�?             @������������������������       �                     @                        ��2>@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @       '                    �?j���� �?             1@       "                     �?      �?             0@                        ��+T@�<ݚ�?             "@������������������������       �                     @        !                   @C@�q�q�?             @������������������������       �                      @������������������������       �                     �?#       &                    �?և���X�?             @$       %                   �7@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?)       �                 `��R@)�n��?�            �v@*       1                    @L�}�:G�?�            `u@+       ,                     @��<b���?             7@������������������������       �        	             0@-       .                 ��A>@����X�?             @������������������������       �                     @/       0                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @2       [                    �?�������?�            �s@3       8                    �?k��9�?3            �V@4       5                    @�eP*L��?             &@������������������������       �                     @6       7                 `f�@      �?              @������������������������       �                     @������������������������       �                     @9       D                     @�����?/            �S@:       C                   �J@ףp=
�?             D@;       <                     �?�}�+r��?             C@������������������������       �                     $@=       >                   �4@@4և���?             <@������������������������       �                     ,@?       @                   @C@؇���X�?	             ,@������������������������       �                     "@A       B                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @E       Z                    �?�(�Tw��?            �C@F       S                    �?
j*D>�?             :@G       R                    <@D�n�3�?             3@H       Q                    �?�n_Y�K�?             *@I       P                 �[$@�q�q�?             (@J       K                 �&B@�<ݚ�?             "@������������������������       �                     @L       M                    0@���Q��?             @������������������������       �                     �?N       O                    3@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @T       Y                 03�9@և���X�?             @U       X                    �?      �?             @V       W                 xFT!@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     *@\       ]                    �?T�����?�            �l@������������������������       �                     6@^       q                 ��) @ƺ"+L�?�            �i@_       p                    �?P��BNֱ?4            �T@`       o                 �?$@���(-�?/            @R@a       b                     @     ��?             @@������������������������       �                      @c       f                 @3�@      �?             8@d       e                    6@      �?              @������������������������       �                     �?������������������������       �                     �?g       h                 ���@�C��2(�?             6@������������������������       �                     @i       j                 ���@�r����?
             .@������������������������       �                     �?k       l                 �|Y=@@4և���?	             ,@������������������������       �                     @m       n                 ���@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �D@������������������������       �                     $@r       s                 pF� @X��Oԣ�?P             _@������������������������       �                     �?t       w                    #@��U!~2�?O            �^@u       v                     @      �?              @������������������������       �                     �?������������������������       �                     �?x       �                    �?�R����?M            @^@y       �                   �<@؇���X�?6             U@z                            @ >�֕�?            �A@{       ~                    4@$�q-�?             :@|       }                    &@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        
             5@������������������������       �                     "@�       �                   �H@�����?"            �H@�       �                 ��1:@      �?             D@�       �                    @@8�Z$���?             :@�       �                   �+@�z�G��?             $@�       �                   �'@���Q��?             @�       �                 �|Y=@�q�q�?             @�       �                    $@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?      �?             0@�       �                     @�8��8��?	             (@�       �                 `fF)@      �?              @������������������������       �                     �?�       �                   @D@؇���X�?             @������������������������       �                     @�       �                   @F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �G@և���X�?	             ,@�       �                   �F@�q�q�?             (@�       �                   �@@      �?              @�       �                   �>@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                    �B@�       �                    @ �q�q�?             8@������������������������       �                     6@�       �                    5@      �?              @������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hR�Bp
       �q@     �c@      ?@     �G@      @      ;@      @      @      �?      @              @      �?               @                      4@      <@      4@      5@      $@      5@       @              @      5@      @      @      @      @              @      @      @                      @      ,@      �?      @      �?      @              �?      �?              �?      �?               @                       @      @      $@      @      $@       @      @              @       @      �?       @                      �?      @      @      @      @              @      @              �?              �?              p@     �[@     �o@     �U@      @      2@              0@      @       @      @              �?       @      �?                       @     @o@     @Q@      C@      J@      @      @      @              @      @              @      @              @@     �G@      @      B@       @      B@              $@       @      :@              ,@       @      (@              "@       @      @       @                      @       @              <@      &@      .@      &@      &@       @      @       @      @      @       @      @              @       @      @      �?              �?      @              @      �?              @                      �?      @              @      @      �?      @      �?       @               @      �?                      �?      @              *@             �j@      1@      6@             �g@      1@      T@      @     �Q@      @      =@      @       @              5@      @      �?      �?      �?                      �?      4@       @      @              *@       @              �?      *@      �?      @              @      �?      @                      �?     �D@              $@             �[@      ,@              �?     �[@      *@      �?      �?      �?                      �?     @[@      (@      R@      (@     �@@       @      8@       @      @       @               @      @              5@              "@             �C@      $@      >@      $@      6@      @      @      @       @      @       @      �?      �?      �?              �?      �?              �?                       @      @              .@      �?      &@      �?      @      �?      �?              @      �?      @              �?      �?              �?      �?              @              @               @      @       @      @      @      @      @      �?              �?      @                      @      @                       @      "@             �B@              �?      7@              6@      �?      �?      �?                      �?r�  tr�  bubhhubehhub.